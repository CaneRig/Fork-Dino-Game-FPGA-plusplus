module bit_stream
(input clk, EA, input [8:0] jump_chn, input [10:0] count_h, count_v, input [11:0] cactuses0, cactuses1, cactuses2, cactuses3, input game_over, output red, blue, green);

reg r = 0;
reg g = 0;
reg b = 0;

integer dino_count;
reg [2:0] dino_sprite_choice = 2;
reg [1:0] dino_sprite [0:3][0:100][0:100];
integer dyno_x, dyno_y;

integer ground_y = 400;

reg [11:0] cactuses [0:4];
integer i = 0;

reg [3:0] cactuses_sprite_choice [0:32];
reg [5:0] choice = 0;
reg [1:0] cactus_sprite [0:7][0:50][0:100];
integer cactus_x, cactus_y;

assign red = r;
assign green = g;
assign blue = b;


always @ (negedge clk)
begin
if (EA) begin

	cactuses[0] = cactuses0;
	cactuses[1] = cactuses1;
	cactuses[2] = cactuses2;
	cactuses[3] = cactuses3;

	if (count_h >= 0) //background
	begin
		r = 0;
		g = 0;
		b = 0;
	end
	
	if (count_v > ground_y-1 & count_v < ground_y + 4) //ground
	begin
		r = 1;
		g = 1;
		b = 1;
	end
		
	dyno_x = count_h - 200;
	dyno_y = 100 - (ground_y - count_v - jump_chn);
  
	// -- DYNO SPRITE --
	dino_sprite[0][2][35] = 1;dino_sprite[0][2][36] = 1;dino_sprite[0][2][37] = 1;dino_sprite[0][2][38] = 1;dino_sprite[0][2][39] = 1;dino_sprite[0][2][40] = 1;dino_sprite[0][2][41] = 1;dino_sprite[0][2][42] = 1;dino_sprite[0][2][43] = 1;dino_sprite[0][2][44] = 1;dino_sprite[0][2][45] = 1;dino_sprite[0][2][46] = 1;dino_sprite[0][2][47] = 1;dino_sprite[0][2][48] = 1;dino_sprite[0][2][49] = 1;dino_sprite[0][2][50] = 1;dino_sprite[0][2][51] = 1;dino_sprite[0][2][52] = 1;dino_sprite[0][2][53] = 1;dino_sprite[0][2][54] = 1;dino_sprite[0][2][55] = 1;dino_sprite[0][2][56] = 1;dino_sprite[0][2][57] = 1;dino_sprite[0][2][58] = 1;dino_sprite[0][2][59] = 1;dino_sprite[0][2][60] = 1;dino_sprite[0][2][61] = 1;dino_sprite[0][2][62] = 1;dino_sprite[0][3][35] = 1;dino_sprite[0][3][36] = 1;dino_sprite[0][3][37] = 1;dino_sprite[0][3][38] = 1;dino_sprite[0][3][39] = 1;dino_sprite[0][3][40] = 1;dino_sprite[0][3][41] = 1;dino_sprite[0][3][42] = 1;dino_sprite[0][3][43] = 1;dino_sprite[0][3][44] = 1;dino_sprite[0][3][45] = 1;dino_sprite[0][3][46] = 1;dino_sprite[0][3][47] = 1;dino_sprite[0][3][48] = 1;dino_sprite[0][3][49] = 1;dino_sprite[0][3][50] = 1;dino_sprite[0][3][51] = 1;dino_sprite[0][3][52] = 1;dino_sprite[0][3][53] = 1;dino_sprite[0][3][54] = 1;dino_sprite[0][3][55] = 1;dino_sprite[0][3][56] = 1;dino_sprite[0][3][57] = 1;dino_sprite[0][3][58] = 1;dino_sprite[0][3][59] = 1;dino_sprite[0][3][60] = 1;dino_sprite[0][3][61] = 1;dino_sprite[0][3][62] = 1;dino_sprite[0][4][35] = 1;dino_sprite[0][4][36] = 1;dino_sprite[0][4][37] = 1;dino_sprite[0][4][38] = 1;dino_sprite[0][4][39] = 1;dino_sprite[0][4][40] = 1;dino_sprite[0][4][41] = 1;dino_sprite[0][4][42] = 1;dino_sprite[0][4][43] = 1;dino_sprite[0][4][44] = 1;dino_sprite[0][4][45] = 1;dino_sprite[0][4][46] = 1;dino_sprite[0][4][47] = 1;dino_sprite[0][4][48] = 1;dino_sprite[0][4][49] = 1;dino_sprite[0][4][50] = 1;dino_sprite[0][4][51] = 1;dino_sprite[0][4][52] = 1;dino_sprite[0][4][53] = 1;dino_sprite[0][4][54] = 1;dino_sprite[0][4][55] = 1;dino_sprite[0][4][56] = 1;dino_sprite[0][4][57] = 1;dino_sprite[0][4][58] = 1;dino_sprite[0][4][59] = 1;dino_sprite[0][4][60] = 1;dino_sprite[0][4][61] = 1;dino_sprite[0][4][62] = 1;dino_sprite[0][5][35] = 1;dino_sprite[0][5][36] = 1;dino_sprite[0][5][37] = 1;dino_sprite[0][5][38] = 1;dino_sprite[0][5][39] = 1;dino_sprite[0][5][40] = 1;dino_sprite[0][5][41] = 1;dino_sprite[0][5][42] = 1;dino_sprite[0][5][43] = 1;dino_sprite[0][5][44] = 1;dino_sprite[0][5][45] = 1;dino_sprite[0][5][46] = 1;dino_sprite[0][5][47] = 1;dino_sprite[0][5][48] = 1;dino_sprite[0][5][49] = 1;dino_sprite[0][5][50] = 1;dino_sprite[0][5][51] = 1;dino_sprite[0][5][52] = 1;dino_sprite[0][5][53] = 1;dino_sprite[0][5][54] = 1;dino_sprite[0][5][55] = 1;dino_sprite[0][5][56] = 1;dino_sprite[0][5][57] = 1;dino_sprite[0][5][58] = 1;dino_sprite[0][5][59] = 1;dino_sprite[0][5][60] = 1;dino_sprite[0][5][61] = 1;dino_sprite[0][5][62] = 1;dino_sprite[0][6][35] = 1;dino_sprite[0][6][36] = 1;dino_sprite[0][6][37] = 1;dino_sprite[0][6][38] = 1;dino_sprite[0][6][39] = 1;dino_sprite[0][6][40] = 1;dino_sprite[0][6][41] = 1;dino_sprite[0][6][42] = 1;dino_sprite[0][6][43] = 1;dino_sprite[0][6][44] = 1;dino_sprite[0][6][45] = 1;dino_sprite[0][6][46] = 1;dino_sprite[0][6][47] = 1;dino_sprite[0][6][48] = 1;dino_sprite[0][6][49] = 1;dino_sprite[0][6][50] = 1;dino_sprite[0][6][51] = 1;dino_sprite[0][6][52] = 1;dino_sprite[0][6][53] = 1;dino_sprite[0][6][54] = 1;dino_sprite[0][6][55] = 1;dino_sprite[0][6][56] = 1;dino_sprite[0][6][57] = 1;dino_sprite[0][6][58] = 1;dino_sprite[0][6][59] = 1;dino_sprite[0][6][60] = 1;dino_sprite[0][6][61] = 1;dino_sprite[0][6][62] = 1;dino_sprite[0][7][35] = 1;dino_sprite[0][7][36] = 1;dino_sprite[0][7][37] = 1;dino_sprite[0][7][38] = 1;dino_sprite[0][7][39] = 1;dino_sprite[0][7][40] = 1;dino_sprite[0][7][41] = 1;dino_sprite[0][7][42] = 1;dino_sprite[0][7][43] = 1;dino_sprite[0][7][44] = 1;dino_sprite[0][7][45] = 1;dino_sprite[0][7][46] = 1;dino_sprite[0][7][47] = 1;dino_sprite[0][7][48] = 1;dino_sprite[0][7][49] = 1;dino_sprite[0][7][50] = 1;dino_sprite[0][7][51] = 1;dino_sprite[0][7][52] = 1;dino_sprite[0][7][53] = 1;dino_sprite[0][7][54] = 1;dino_sprite[0][7][55] = 1;dino_sprite[0][7][56] = 1;dino_sprite[0][7][57] = 1;dino_sprite[0][7][58] = 1;dino_sprite[0][7][59] = 1;dino_sprite[0][7][60] = 1;dino_sprite[0][7][61] = 1;dino_sprite[0][7][62] = 1;dino_sprite[0][7][63] = 1;dino_sprite[0][7][64] = 1;dino_sprite[0][7][65] = 1;dino_sprite[0][7][66] = 1;dino_sprite[0][7][67] = 1;dino_sprite[0][8][44] = 1;dino_sprite[0][8][45] = 1;dino_sprite[0][8][46] = 1;dino_sprite[0][8][47] = 1;dino_sprite[0][8][48] = 1;dino_sprite[0][8][49] = 1;dino_sprite[0][8][50] = 1;dino_sprite[0][8][51] = 1;dino_sprite[0][8][52] = 1;dino_sprite[0][8][53] = 1;dino_sprite[0][8][54] = 1;dino_sprite[0][8][55] = 1;dino_sprite[0][8][56] = 1;dino_sprite[0][8][57] = 1;dino_sprite[0][8][58] = 1;dino_sprite[0][8][59] = 1;dino_sprite[0][8][60] = 1;dino_sprite[0][8][61] = 1;dino_sprite[0][8][62] = 1;dino_sprite[0][8][63] = 1;dino_sprite[0][8][64] = 1;dino_sprite[0][8][65] = 1;dino_sprite[0][8][66] = 1;dino_sprite[0][8][67] = 1;dino_sprite[0][9][44] = 1;dino_sprite[0][9][45] = 1;dino_sprite[0][9][46] = 1;dino_sprite[0][9][47] = 1;dino_sprite[0][9][48] = 1;dino_sprite[0][9][49] = 1;dino_sprite[0][9][50] = 1;dino_sprite[0][9][51] = 1;dino_sprite[0][9][52] = 1;dino_sprite[0][9][53] = 1;dino_sprite[0][9][54] = 1;dino_sprite[0][9][55] = 1;dino_sprite[0][9][56] = 1;dino_sprite[0][9][57] = 1;dino_sprite[0][9][58] = 1;dino_sprite[0][9][59] = 1;dino_sprite[0][9][60] = 1;dino_sprite[0][9][61] = 1;dino_sprite[0][9][62] = 1;dino_sprite[0][9][63] = 1;dino_sprite[0][9][64] = 1;dino_sprite[0][9][65] = 1;dino_sprite[0][9][66] = 1;dino_sprite[0][9][67] = 1;dino_sprite[0][10][44] = 1;dino_sprite[0][10][45] = 1;dino_sprite[0][10][46] = 1;dino_sprite[0][10][47] = 1;dino_sprite[0][10][48] = 1;dino_sprite[0][10][49] = 1;dino_sprite[0][10][50] = 1;dino_sprite[0][10][51] = 1;dino_sprite[0][10][52] = 1;dino_sprite[0][10][53] = 1;dino_sprite[0][10][54] = 1;dino_sprite[0][10][55] = 1;dino_sprite[0][10][56] = 1;dino_sprite[0][10][57] = 1;dino_sprite[0][10][58] = 1;dino_sprite[0][10][59] = 1;dino_sprite[0][10][60] = 1;dino_sprite[0][10][61] = 1;dino_sprite[0][10][62] = 1;dino_sprite[0][10][63] = 1;dino_sprite[0][10][64] = 1;dino_sprite[0][10][65] = 1;dino_sprite[0][10][66] = 1;dino_sprite[0][10][67] = 1;dino_sprite[0][11][44] = 1;dino_sprite[0][11][45] = 1;dino_sprite[0][11][46] = 1;dino_sprite[0][11][47] = 1;dino_sprite[0][11][48] = 1;dino_sprite[0][11][49] = 1;dino_sprite[0][11][50] = 1;dino_sprite[0][11][51] = 1;dino_sprite[0][11][52] = 1;dino_sprite[0][11][53] = 1;dino_sprite[0][11][54] = 1;dino_sprite[0][11][55] = 1;dino_sprite[0][11][56] = 1;dino_sprite[0][11][57] = 1;dino_sprite[0][11][58] = 1;dino_sprite[0][11][59] = 1;dino_sprite[0][11][60] = 1;dino_sprite[0][11][61] = 1;dino_sprite[0][11][62] = 1;dino_sprite[0][11][63] = 1;dino_sprite[0][11][64] = 1;dino_sprite[0][11][65] = 1;dino_sprite[0][11][66] = 1;dino_sprite[0][11][67] = 1;dino_sprite[0][12][49] = 1;dino_sprite[0][12][50] = 1;dino_sprite[0][12][51] = 1;dino_sprite[0][12][52] = 1;dino_sprite[0][12][53] = 1;dino_sprite[0][12][54] = 1;dino_sprite[0][12][55] = 1;dino_sprite[0][12][56] = 1;dino_sprite[0][12][57] = 1;dino_sprite[0][12][58] = 1;dino_sprite[0][12][59] = 1;dino_sprite[0][12][60] = 1;dino_sprite[0][12][61] = 1;dino_sprite[0][12][62] = 1;dino_sprite[0][12][63] = 1;dino_sprite[0][12][64] = 1;dino_sprite[0][12][65] = 1;dino_sprite[0][12][66] = 1;dino_sprite[0][12][67] = 1;dino_sprite[0][12][68] = 1;dino_sprite[0][12][69] = 1;dino_sprite[0][12][70] = 1;dino_sprite[0][12][71] = 1;dino_sprite[0][12][72] = 1;dino_sprite[0][13][49] = 1;dino_sprite[0][13][50] = 1;dino_sprite[0][13][51] = 1;dino_sprite[0][13][52] = 1;dino_sprite[0][13][53] = 1;dino_sprite[0][13][54] = 1;dino_sprite[0][13][55] = 1;dino_sprite[0][13][56] = 1;dino_sprite[0][13][57] = 1;dino_sprite[0][13][58] = 1;dino_sprite[0][13][59] = 1;dino_sprite[0][13][60] = 1;dino_sprite[0][13][61] = 1;dino_sprite[0][13][62] = 1;dino_sprite[0][13][63] = 1;dino_sprite[0][13][64] = 1;dino_sprite[0][13][65] = 1;dino_sprite[0][13][66] = 1;dino_sprite[0][13][67] = 1;dino_sprite[0][13][68] = 1;dino_sprite[0][13][69] = 1;dino_sprite[0][13][70] = 1;dino_sprite[0][13][71] = 1;dino_sprite[0][13][72] = 1;dino_sprite[0][14][49] = 1;dino_sprite[0][14][50] = 1;dino_sprite[0][14][51] = 1;dino_sprite[0][14][52] = 1;dino_sprite[0][14][53] = 1;dino_sprite[0][14][54] = 1;dino_sprite[0][14][55] = 1;dino_sprite[0][14][56] = 1;dino_sprite[0][14][57] = 1;dino_sprite[0][14][58] = 1;dino_sprite[0][14][59] = 1;dino_sprite[0][14][60] = 1;dino_sprite[0][14][61] = 1;dino_sprite[0][14][62] = 1;dino_sprite[0][14][63] = 1;dino_sprite[0][14][64] = 1;dino_sprite[0][14][65] = 1;dino_sprite[0][14][66] = 1;dino_sprite[0][14][67] = 1;dino_sprite[0][14][68] = 1;dino_sprite[0][14][69] = 1;dino_sprite[0][14][70] = 1;dino_sprite[0][14][71] = 1;dino_sprite[0][14][72] = 1;dino_sprite[0][15][49] = 1;dino_sprite[0][15][50] = 1;dino_sprite[0][15][51] = 1;dino_sprite[0][15][52] = 1;dino_sprite[0][15][53] = 1;dino_sprite[0][15][54] = 1;dino_sprite[0][15][55] = 1;dino_sprite[0][15][56] = 1;dino_sprite[0][15][57] = 1;dino_sprite[0][15][58] = 1;dino_sprite[0][15][59] = 1;dino_sprite[0][15][60] = 1;dino_sprite[0][15][61] = 1;dino_sprite[0][15][62] = 1;dino_sprite[0][15][63] = 1;dino_sprite[0][15][64] = 1;dino_sprite[0][15][65] = 1;dino_sprite[0][15][66] = 1;dino_sprite[0][15][67] = 1;dino_sprite[0][15][68] = 1;dino_sprite[0][15][69] = 1;dino_sprite[0][15][70] = 1;dino_sprite[0][15][71] = 1;dino_sprite[0][15][72] = 1;dino_sprite[0][16][49] = 1;dino_sprite[0][16][50] = 1;dino_sprite[0][16][51] = 1;dino_sprite[0][16][52] = 1;dino_sprite[0][16][53] = 1;dino_sprite[0][16][54] = 1;dino_sprite[0][16][55] = 1;dino_sprite[0][16][56] = 1;dino_sprite[0][16][57] = 1;dino_sprite[0][16][58] = 1;dino_sprite[0][16][59] = 1;dino_sprite[0][16][60] = 1;dino_sprite[0][16][61] = 1;dino_sprite[0][16][62] = 1;dino_sprite[0][16][63] = 1;dino_sprite[0][16][64] = 1;dino_sprite[0][16][65] = 1;dino_sprite[0][16][66] = 1;dino_sprite[0][16][67] = 1;dino_sprite[0][16][68] = 1;dino_sprite[0][16][69] = 1;dino_sprite[0][16][70] = 1;dino_sprite[0][16][71] = 1;dino_sprite[0][16][72] = 1;dino_sprite[0][17][54] = 1;dino_sprite[0][17][55] = 1;dino_sprite[0][17][56] = 1;dino_sprite[0][17][57] = 1;dino_sprite[0][17][58] = 1;dino_sprite[0][17][59] = 1;dino_sprite[0][17][60] = 1;dino_sprite[0][17][61] = 1;dino_sprite[0][17][62] = 1;dino_sprite[0][17][63] = 1;dino_sprite[0][17][64] = 1;dino_sprite[0][17][65] = 1;dino_sprite[0][17][66] = 1;dino_sprite[0][17][67] = 1;dino_sprite[0][17][68] = 1;dino_sprite[0][17][69] = 1;dino_sprite[0][17][70] = 1;dino_sprite[0][17][71] = 1;dino_sprite[0][17][72] = 1;dino_sprite[0][17][73] = 1;dino_sprite[0][17][74] = 1;dino_sprite[0][17][75] = 1;dino_sprite[0][17][76] = 1;dino_sprite[0][17][77] = 1;dino_sprite[0][18][54] = 1;dino_sprite[0][18][55] = 1;dino_sprite[0][18][56] = 1;dino_sprite[0][18][57] = 1;dino_sprite[0][18][58] = 1;dino_sprite[0][18][59] = 1;dino_sprite[0][18][60] = 1;dino_sprite[0][18][61] = 1;dino_sprite[0][18][62] = 1;dino_sprite[0][18][63] = 1;dino_sprite[0][18][64] = 1;dino_sprite[0][18][65] = 1;dino_sprite[0][18][66] = 1;dino_sprite[0][18][67] = 1;dino_sprite[0][18][68] = 1;dino_sprite[0][18][69] = 1;dino_sprite[0][18][70] = 1;dino_sprite[0][18][71] = 1;dino_sprite[0][18][72] = 1;dino_sprite[0][18][73] = 1;dino_sprite[0][18][74] = 1;dino_sprite[0][18][75] = 1;dino_sprite[0][18][76] = 1;dino_sprite[0][18][77] = 1;dino_sprite[0][19][54] = 1;dino_sprite[0][19][55] = 1;dino_sprite[0][19][56] = 1;dino_sprite[0][19][57] = 1;dino_sprite[0][19][58] = 1;dino_sprite[0][19][59] = 1;dino_sprite[0][19][60] = 1;dino_sprite[0][19][61] = 1;dino_sprite[0][19][62] = 1;dino_sprite[0][19][63] = 1;dino_sprite[0][19][64] = 1;dino_sprite[0][19][65] = 1;dino_sprite[0][19][66] = 1;dino_sprite[0][19][67] = 1;dino_sprite[0][19][68] = 1;dino_sprite[0][19][69] = 1;dino_sprite[0][19][70] = 1;dino_sprite[0][19][71] = 1;dino_sprite[0][19][72] = 1;dino_sprite[0][19][73] = 1;dino_sprite[0][19][74] = 1;dino_sprite[0][19][75] = 1;dino_sprite[0][19][76] = 1;dino_sprite[0][19][77] = 1;dino_sprite[0][20][54] = 1;dino_sprite[0][20][55] = 1;dino_sprite[0][20][56] = 1;dino_sprite[0][20][57] = 1;dino_sprite[0][20][58] = 1;dino_sprite[0][20][59] = 1;dino_sprite[0][20][60] = 1;dino_sprite[0][20][61] = 1;dino_sprite[0][20][62] = 1;dino_sprite[0][20][63] = 1;dino_sprite[0][20][64] = 1;dino_sprite[0][20][65] = 1;dino_sprite[0][20][66] = 1;dino_sprite[0][20][67] = 1;dino_sprite[0][20][68] = 1;dino_sprite[0][20][69] = 1;dino_sprite[0][20][70] = 1;dino_sprite[0][20][71] = 1;dino_sprite[0][20][72] = 1;dino_sprite[0][20][73] = 1;dino_sprite[0][20][74] = 1;dino_sprite[0][20][75] = 1;dino_sprite[0][20][76] = 1;dino_sprite[0][20][77] = 1;dino_sprite[0][21][54] = 1;dino_sprite[0][21][55] = 1;dino_sprite[0][21][56] = 1;dino_sprite[0][21][57] = 1;dino_sprite[0][21][58] = 1;dino_sprite[0][21][59] = 1;dino_sprite[0][21][60] = 1;dino_sprite[0][21][61] = 1;dino_sprite[0][21][62] = 1;dino_sprite[0][21][63] = 1;dino_sprite[0][21][64] = 1;dino_sprite[0][21][65] = 1;dino_sprite[0][21][66] = 1;dino_sprite[0][21][67] = 1;dino_sprite[0][21][68] = 1;dino_sprite[0][21][69] = 1;dino_sprite[0][21][70] = 1;dino_sprite[0][21][71] = 1;dino_sprite[0][21][72] = 1;dino_sprite[0][21][73] = 1;dino_sprite[0][21][74] = 1;dino_sprite[0][21][75] = 1;dino_sprite[0][21][76] = 1;dino_sprite[0][21][77] = 1;dino_sprite[0][22][54] = 1;dino_sprite[0][22][55] = 1;dino_sprite[0][22][56] = 1;dino_sprite[0][22][57] = 1;dino_sprite[0][22][58] = 1;dino_sprite[0][22][59] = 1;dino_sprite[0][22][60] = 1;dino_sprite[0][22][61] = 1;dino_sprite[0][22][62] = 1;dino_sprite[0][22][63] = 1;dino_sprite[0][22][64] = 1;dino_sprite[0][22][65] = 1;dino_sprite[0][22][66] = 1;dino_sprite[0][22][67] = 1;dino_sprite[0][22][68] = 1;dino_sprite[0][22][69] = 1;dino_sprite[0][22][70] = 1;dino_sprite[0][22][71] = 1;dino_sprite[0][22][72] = 1;dino_sprite[0][22][73] = 1;dino_sprite[0][22][74] = 1;dino_sprite[0][22][75] = 1;dino_sprite[0][22][76] = 1;dino_sprite[0][22][77] = 1;dino_sprite[0][22][78] = 1;dino_sprite[0][22][79] = 1;dino_sprite[0][22][80] = 1;dino_sprite[0][22][81] = 1;dino_sprite[0][23][54] = 1;dino_sprite[0][23][55] = 1;dino_sprite[0][23][56] = 1;dino_sprite[0][23][57] = 1;dino_sprite[0][23][58] = 1;dino_sprite[0][23][59] = 1;dino_sprite[0][23][60] = 1;dino_sprite[0][23][61] = 1;dino_sprite[0][23][62] = 1;dino_sprite[0][23][63] = 1;dino_sprite[0][23][64] = 1;dino_sprite[0][23][65] = 1;dino_sprite[0][23][66] = 1;dino_sprite[0][23][67] = 1;dino_sprite[0][23][68] = 1;dino_sprite[0][23][69] = 1;dino_sprite[0][23][70] = 1;dino_sprite[0][23][71] = 1;dino_sprite[0][23][72] = 1;dino_sprite[0][23][73] = 1;dino_sprite[0][23][74] = 1;dino_sprite[0][23][75] = 1;dino_sprite[0][23][76] = 1;dino_sprite[0][23][77] = 1;dino_sprite[0][23][78] = 1;dino_sprite[0][23][79] = 1;dino_sprite[0][23][80] = 1;dino_sprite[0][23][81] = 1;dino_sprite[0][24][54] = 1;dino_sprite[0][24][55] = 1;dino_sprite[0][24][56] = 1;dino_sprite[0][24][57] = 1;dino_sprite[0][24][58] = 1;dino_sprite[0][24][59] = 1;dino_sprite[0][24][60] = 1;dino_sprite[0][24][61] = 1;dino_sprite[0][24][62] = 1;dino_sprite[0][24][63] = 1;dino_sprite[0][24][64] = 1;dino_sprite[0][24][65] = 1;dino_sprite[0][24][66] = 1;dino_sprite[0][24][67] = 1;dino_sprite[0][24][68] = 1;dino_sprite[0][24][69] = 1;dino_sprite[0][24][70] = 1;dino_sprite[0][24][71] = 1;dino_sprite[0][24][72] = 1;dino_sprite[0][24][73] = 1;dino_sprite[0][24][74] = 1;dino_sprite[0][24][75] = 1;dino_sprite[0][24][76] = 1;dino_sprite[0][24][77] = 1;dino_sprite[0][24][78] = 1;dino_sprite[0][24][79] = 1;dino_sprite[0][24][80] = 1;dino_sprite[0][24][81] = 1;dino_sprite[0][25][54] = 1;dino_sprite[0][25][55] = 1;dino_sprite[0][25][56] = 1;dino_sprite[0][25][57] = 1;dino_sprite[0][25][58] = 1;dino_sprite[0][25][59] = 1;dino_sprite[0][25][60] = 1;dino_sprite[0][25][61] = 1;dino_sprite[0][25][62] = 1;dino_sprite[0][25][63] = 1;dino_sprite[0][25][64] = 1;dino_sprite[0][25][65] = 1;dino_sprite[0][25][66] = 1;dino_sprite[0][25][67] = 1;dino_sprite[0][25][68] = 1;dino_sprite[0][25][69] = 1;dino_sprite[0][25][70] = 1;dino_sprite[0][25][71] = 1;dino_sprite[0][25][72] = 1;dino_sprite[0][25][73] = 1;dino_sprite[0][25][74] = 1;dino_sprite[0][25][75] = 1;dino_sprite[0][25][76] = 1;dino_sprite[0][25][77] = 1;dino_sprite[0][25][78] = 1;dino_sprite[0][25][79] = 1;dino_sprite[0][25][80] = 1;dino_sprite[0][25][81] = 1;dino_sprite[0][26][49] = 1;dino_sprite[0][26][50] = 1;dino_sprite[0][26][51] = 1;dino_sprite[0][26][52] = 1;dino_sprite[0][26][53] = 1;dino_sprite[0][26][54] = 1;dino_sprite[0][26][55] = 1;dino_sprite[0][26][56] = 1;dino_sprite[0][26][57] = 1;dino_sprite[0][26][58] = 1;dino_sprite[0][26][59] = 1;dino_sprite[0][26][60] = 1;dino_sprite[0][26][61] = 1;dino_sprite[0][26][62] = 1;dino_sprite[0][26][63] = 1;dino_sprite[0][26][64] = 1;dino_sprite[0][26][65] = 1;dino_sprite[0][26][66] = 1;dino_sprite[0][26][67] = 1;dino_sprite[0][26][68] = 1;dino_sprite[0][26][69] = 1;dino_sprite[0][26][70] = 1;dino_sprite[0][26][71] = 1;dino_sprite[0][26][72] = 1;dino_sprite[0][26][73] = 1;dino_sprite[0][26][74] = 1;dino_sprite[0][26][75] = 1;dino_sprite[0][26][76] = 1;dino_sprite[0][26][77] = 1;dino_sprite[0][26][78] = 1;dino_sprite[0][26][79] = 1;dino_sprite[0][26][80] = 1;dino_sprite[0][26][81] = 1;dino_sprite[0][26][82] = 1;dino_sprite[0][26][83] = 1;dino_sprite[0][26][84] = 1;dino_sprite[0][26][85] = 1;dino_sprite[0][26][86] = 1;dino_sprite[0][26][87] = 1;dino_sprite[0][26][88] = 1;dino_sprite[0][26][89] = 1;dino_sprite[0][26][90] = 1;dino_sprite[0][26][91] = 1;dino_sprite[0][26][92] = 1;dino_sprite[0][26][93] = 1;dino_sprite[0][26][94] = 1;dino_sprite[0][26][95] = 1;dino_sprite[0][26][96] = 1;dino_sprite[0][26][97] = 1;dino_sprite[0][26][98] = 1;dino_sprite[0][26][99] = 1;dino_sprite[0][27][49] = 1;dino_sprite[0][27][50] = 1;dino_sprite[0][27][51] = 1;dino_sprite[0][27][52] = 1;dino_sprite[0][27][53] = 1;dino_sprite[0][27][54] = 1;dino_sprite[0][27][55] = 1;dino_sprite[0][27][56] = 1;dino_sprite[0][27][57] = 1;dino_sprite[0][27][58] = 1;dino_sprite[0][27][59] = 1;dino_sprite[0][27][60] = 1;dino_sprite[0][27][61] = 1;dino_sprite[0][27][62] = 1;dino_sprite[0][27][63] = 1;dino_sprite[0][27][64] = 1;dino_sprite[0][27][65] = 1;dino_sprite[0][27][66] = 1;dino_sprite[0][27][67] = 1;dino_sprite[0][27][68] = 1;dino_sprite[0][27][69] = 1;dino_sprite[0][27][70] = 1;dino_sprite[0][27][71] = 1;dino_sprite[0][27][72] = 1;dino_sprite[0][27][73] = 1;dino_sprite[0][27][74] = 1;dino_sprite[0][27][75] = 1;dino_sprite[0][27][76] = 1;dino_sprite[0][27][77] = 1;dino_sprite[0][27][78] = 1;dino_sprite[0][27][79] = 1;dino_sprite[0][27][80] = 1;dino_sprite[0][27][81] = 1;dino_sprite[0][27][82] = 1;dino_sprite[0][27][83] = 1;dino_sprite[0][27][84] = 1;dino_sprite[0][27][85] = 1;dino_sprite[0][27][86] = 1;dino_sprite[0][27][87] = 1;dino_sprite[0][27][88] = 1;dino_sprite[0][27][89] = 1;dino_sprite[0][27][90] = 1;dino_sprite[0][27][91] = 1;dino_sprite[0][27][92] = 1;dino_sprite[0][27][93] = 1;dino_sprite[0][27][94] = 1;dino_sprite[0][27][95] = 1;dino_sprite[0][27][96] = 1;dino_sprite[0][27][97] = 1;dino_sprite[0][27][98] = 1;dino_sprite[0][27][99] = 1;dino_sprite[0][28][49] = 1;dino_sprite[0][28][50] = 1;dino_sprite[0][28][51] = 1;dino_sprite[0][28][52] = 1;dino_sprite[0][28][53] = 1;dino_sprite[0][28][54] = 1;dino_sprite[0][28][55] = 1;dino_sprite[0][28][56] = 1;dino_sprite[0][28][57] = 1;dino_sprite[0][28][58] = 1;dino_sprite[0][28][59] = 1;dino_sprite[0][28][60] = 1;dino_sprite[0][28][61] = 1;dino_sprite[0][28][62] = 1;dino_sprite[0][28][63] = 1;dino_sprite[0][28][64] = 1;dino_sprite[0][28][65] = 1;dino_sprite[0][28][66] = 1;dino_sprite[0][28][67] = 1;dino_sprite[0][28][68] = 1;dino_sprite[0][28][69] = 1;dino_sprite[0][28][70] = 1;dino_sprite[0][28][71] = 1;dino_sprite[0][28][72] = 1;dino_sprite[0][28][73] = 1;dino_sprite[0][28][74] = 1;dino_sprite[0][28][75] = 1;dino_sprite[0][28][76] = 1;dino_sprite[0][28][77] = 1;dino_sprite[0][28][78] = 1;dino_sprite[0][28][79] = 1;dino_sprite[0][28][80] = 1;dino_sprite[0][28][81] = 1;dino_sprite[0][28][82] = 1;dino_sprite[0][28][83] = 1;dino_sprite[0][28][84] = 1;dino_sprite[0][28][85] = 1;dino_sprite[0][28][86] = 1;dino_sprite[0][28][87] = 1;dino_sprite[0][28][88] = 1;dino_sprite[0][28][89] = 1;dino_sprite[0][28][90] = 1;dino_sprite[0][28][91] = 1;dino_sprite[0][28][92] = 1;dino_sprite[0][28][93] = 1;dino_sprite[0][28][94] = 1;dino_sprite[0][28][95] = 1;dino_sprite[0][28][96] = 1;dino_sprite[0][28][97] = 1;dino_sprite[0][28][98] = 1;dino_sprite[0][28][99] = 1;dino_sprite[0][29][49] = 1;dino_sprite[0][29][50] = 1;dino_sprite[0][29][51] = 1;dino_sprite[0][29][52] = 1;dino_sprite[0][29][53] = 1;dino_sprite[0][29][54] = 1;dino_sprite[0][29][55] = 1;dino_sprite[0][29][56] = 1;dino_sprite[0][29][57] = 1;dino_sprite[0][29][58] = 1;dino_sprite[0][29][59] = 1;dino_sprite[0][29][60] = 1;dino_sprite[0][29][61] = 1;dino_sprite[0][29][62] = 1;dino_sprite[0][29][63] = 1;dino_sprite[0][29][64] = 1;dino_sprite[0][29][65] = 1;dino_sprite[0][29][66] = 1;dino_sprite[0][29][67] = 1;dino_sprite[0][29][68] = 1;dino_sprite[0][29][69] = 1;dino_sprite[0][29][70] = 1;dino_sprite[0][29][71] = 1;dino_sprite[0][29][72] = 1;dino_sprite[0][29][73] = 1;dino_sprite[0][29][74] = 1;dino_sprite[0][29][75] = 1;dino_sprite[0][29][76] = 1;dino_sprite[0][29][77] = 1;dino_sprite[0][29][78] = 1;dino_sprite[0][29][79] = 1;dino_sprite[0][29][80] = 1;dino_sprite[0][29][81] = 1;dino_sprite[0][29][82] = 1;dino_sprite[0][29][83] = 1;dino_sprite[0][29][84] = 1;dino_sprite[0][29][85] = 1;dino_sprite[0][29][86] = 1;dino_sprite[0][29][87] = 1;dino_sprite[0][29][88] = 1;dino_sprite[0][29][89] = 1;dino_sprite[0][29][90] = 1;dino_sprite[0][29][91] = 1;dino_sprite[0][29][92] = 1;dino_sprite[0][29][93] = 1;dino_sprite[0][29][94] = 1;dino_sprite[0][29][95] = 1;dino_sprite[0][29][96] = 1;dino_sprite[0][29][97] = 1;dino_sprite[0][29][98] = 1;dino_sprite[0][29][99] = 1;dino_sprite[0][30][49] = 1;dino_sprite[0][30][50] = 1;dino_sprite[0][30][51] = 1;dino_sprite[0][30][52] = 1;dino_sprite[0][30][53] = 1;dino_sprite[0][30][54] = 1;dino_sprite[0][30][55] = 1;dino_sprite[0][30][56] = 1;dino_sprite[0][30][57] = 1;dino_sprite[0][30][58] = 1;dino_sprite[0][30][59] = 1;dino_sprite[0][30][60] = 1;dino_sprite[0][30][61] = 1;dino_sprite[0][30][62] = 1;dino_sprite[0][30][63] = 1;dino_sprite[0][30][64] = 1;dino_sprite[0][30][65] = 1;dino_sprite[0][30][66] = 1;dino_sprite[0][30][67] = 1;dino_sprite[0][30][68] = 1;dino_sprite[0][30][69] = 1;dino_sprite[0][30][70] = 1;dino_sprite[0][30][71] = 1;dino_sprite[0][30][72] = 1;dino_sprite[0][30][73] = 1;dino_sprite[0][30][74] = 1;dino_sprite[0][30][75] = 1;dino_sprite[0][30][76] = 1;dino_sprite[0][30][77] = 1;dino_sprite[0][30][78] = 1;dino_sprite[0][30][79] = 1;dino_sprite[0][30][80] = 1;dino_sprite[0][30][81] = 1;dino_sprite[0][30][82] = 1;dino_sprite[0][30][83] = 1;dino_sprite[0][30][84] = 1;dino_sprite[0][30][85] = 1;dino_sprite[0][30][86] = 1;dino_sprite[0][30][87] = 1;dino_sprite[0][30][88] = 1;dino_sprite[0][30][89] = 1;dino_sprite[0][30][90] = 1;dino_sprite[0][30][91] = 1;dino_sprite[0][30][92] = 1;dino_sprite[0][30][93] = 1;dino_sprite[0][30][94] = 1;dino_sprite[0][30][95] = 1;dino_sprite[0][30][96] = 1;dino_sprite[0][30][97] = 1;dino_sprite[0][30][98] = 1;dino_sprite[0][30][99] = 1;dino_sprite[0][31][44] = 1;dino_sprite[0][31][45] = 1;dino_sprite[0][31][46] = 1;dino_sprite[0][31][47] = 1;dino_sprite[0][31][48] = 1;dino_sprite[0][31][49] = 1;dino_sprite[0][31][50] = 1;dino_sprite[0][31][51] = 1;dino_sprite[0][31][52] = 1;dino_sprite[0][31][53] = 1;dino_sprite[0][31][54] = 1;dino_sprite[0][31][55] = 1;dino_sprite[0][31][56] = 1;dino_sprite[0][31][57] = 1;dino_sprite[0][31][58] = 1;dino_sprite[0][31][59] = 1;dino_sprite[0][31][60] = 1;dino_sprite[0][31][61] = 1;dino_sprite[0][31][62] = 1;dino_sprite[0][31][63] = 1;dino_sprite[0][31][64] = 1;dino_sprite[0][31][65] = 1;dino_sprite[0][31][66] = 1;dino_sprite[0][31][67] = 1;dino_sprite[0][31][68] = 1;dino_sprite[0][31][69] = 1;dino_sprite[0][31][70] = 1;dino_sprite[0][31][71] = 1;dino_sprite[0][31][72] = 1;dino_sprite[0][31][73] = 1;dino_sprite[0][31][74] = 1;dino_sprite[0][31][75] = 1;dino_sprite[0][31][76] = 1;dino_sprite[0][31][77] = 1;dino_sprite[0][31][78] = 1;dino_sprite[0][31][79] = 1;dino_sprite[0][31][80] = 1;dino_sprite[0][31][81] = 1;dino_sprite[0][31][82] = 1;dino_sprite[0][31][83] = 1;dino_sprite[0][31][84] = 1;dino_sprite[0][31][85] = 1;dino_sprite[0][31][86] = 1;dino_sprite[0][31][87] = 1;dino_sprite[0][31][88] = 1;dino_sprite[0][31][89] = 1;dino_sprite[0][31][90] = 1;dino_sprite[0][31][91] = 1;dino_sprite[0][31][92] = 1;dino_sprite[0][31][93] = 1;dino_sprite[0][31][94] = 1;dino_sprite[0][31][95] = 1;dino_sprite[0][31][96] = 1;dino_sprite[0][31][97] = 1;dino_sprite[0][31][98] = 1;dino_sprite[0][31][99] = 1;dino_sprite[0][32][44] = 1;dino_sprite[0][32][45] = 1;dino_sprite[0][32][46] = 1;dino_sprite[0][32][47] = 1;dino_sprite[0][32][48] = 1;dino_sprite[0][32][49] = 1;dino_sprite[0][32][50] = 1;dino_sprite[0][32][51] = 1;dino_sprite[0][32][52] = 1;dino_sprite[0][32][53] = 1;dino_sprite[0][32][54] = 1;dino_sprite[0][32][55] = 1;dino_sprite[0][32][56] = 1;dino_sprite[0][32][57] = 1;dino_sprite[0][32][58] = 1;dino_sprite[0][32][59] = 1;dino_sprite[0][32][60] = 1;dino_sprite[0][32][61] = 1;dino_sprite[0][32][62] = 1;dino_sprite[0][32][63] = 1;dino_sprite[0][32][64] = 1;dino_sprite[0][32][65] = 1;dino_sprite[0][32][66] = 1;dino_sprite[0][32][67] = 1;dino_sprite[0][32][68] = 1;dino_sprite[0][32][69] = 1;dino_sprite[0][32][70] = 1;dino_sprite[0][32][71] = 1;dino_sprite[0][32][72] = 1;dino_sprite[0][32][73] = 1;dino_sprite[0][32][74] = 1;dino_sprite[0][32][75] = 1;dino_sprite[0][32][76] = 1;dino_sprite[0][32][77] = 1;dino_sprite[0][32][78] = 1;dino_sprite[0][32][79] = 1;dino_sprite[0][32][80] = 1;dino_sprite[0][32][81] = 1;dino_sprite[0][32][82] = 1;dino_sprite[0][32][83] = 1;dino_sprite[0][32][84] = 1;dino_sprite[0][32][85] = 1;dino_sprite[0][32][86] = 1;dino_sprite[0][32][95] = 1;dino_sprite[0][32][96] = 1;dino_sprite[0][32][97] = 1;dino_sprite[0][32][98] = 1;dino_sprite[0][32][99] = 1;dino_sprite[0][33][44] = 1;dino_sprite[0][33][45] = 1;dino_sprite[0][33][46] = 1;dino_sprite[0][33][47] = 1;dino_sprite[0][33][48] = 1;dino_sprite[0][33][49] = 1;dino_sprite[0][33][50] = 1;dino_sprite[0][33][51] = 1;dino_sprite[0][33][52] = 1;dino_sprite[0][33][53] = 1;dino_sprite[0][33][54] = 1;dino_sprite[0][33][55] = 1;dino_sprite[0][33][56] = 1;dino_sprite[0][33][57] = 1;dino_sprite[0][33][58] = 1;dino_sprite[0][33][59] = 1;dino_sprite[0][33][60] = 1;dino_sprite[0][33][61] = 1;dino_sprite[0][33][62] = 1;dino_sprite[0][33][63] = 1;dino_sprite[0][33][64] = 1;dino_sprite[0][33][65] = 1;dino_sprite[0][33][66] = 1;dino_sprite[0][33][67] = 1;dino_sprite[0][33][68] = 1;dino_sprite[0][33][69] = 1;dino_sprite[0][33][70] = 1;dino_sprite[0][33][71] = 1;dino_sprite[0][33][72] = 1;dino_sprite[0][33][73] = 1;dino_sprite[0][33][74] = 1;dino_sprite[0][33][75] = 1;dino_sprite[0][33][76] = 1;dino_sprite[0][33][77] = 1;dino_sprite[0][33][78] = 1;dino_sprite[0][33][79] = 1;dino_sprite[0][33][80] = 1;dino_sprite[0][33][81] = 1;dino_sprite[0][33][82] = 1;dino_sprite[0][33][83] = 1;dino_sprite[0][33][84] = 1;dino_sprite[0][33][85] = 1;dino_sprite[0][33][86] = 1;dino_sprite[0][33][95] = 1;dino_sprite[0][33][96] = 1;dino_sprite[0][33][97] = 1;dino_sprite[0][33][98] = 1;dino_sprite[0][33][99] = 1;dino_sprite[0][34][44] = 1;dino_sprite[0][34][45] = 1;dino_sprite[0][34][46] = 1;dino_sprite[0][34][47] = 1;dino_sprite[0][34][48] = 1;dino_sprite[0][34][49] = 1;dino_sprite[0][34][50] = 1;dino_sprite[0][34][51] = 1;dino_sprite[0][34][52] = 1;dino_sprite[0][34][53] = 1;dino_sprite[0][34][54] = 1;dino_sprite[0][34][55] = 1;dino_sprite[0][34][56] = 1;dino_sprite[0][34][57] = 1;dino_sprite[0][34][58] = 1;dino_sprite[0][34][59] = 1;dino_sprite[0][34][60] = 1;dino_sprite[0][34][61] = 1;dino_sprite[0][34][62] = 1;dino_sprite[0][34][63] = 1;dino_sprite[0][34][64] = 1;dino_sprite[0][34][65] = 1;dino_sprite[0][34][66] = 1;dino_sprite[0][34][67] = 1;dino_sprite[0][34][68] = 1;dino_sprite[0][34][69] = 1;dino_sprite[0][34][70] = 1;dino_sprite[0][34][71] = 1;dino_sprite[0][34][72] = 1;dino_sprite[0][34][73] = 1;dino_sprite[0][34][74] = 1;dino_sprite[0][34][75] = 1;dino_sprite[0][34][76] = 1;dino_sprite[0][34][77] = 1;dino_sprite[0][34][78] = 1;dino_sprite[0][34][79] = 1;dino_sprite[0][34][80] = 1;dino_sprite[0][34][81] = 1;dino_sprite[0][34][82] = 1;dino_sprite[0][34][83] = 1;dino_sprite[0][34][84] = 1;dino_sprite[0][34][85] = 1;dino_sprite[0][34][86] = 1;dino_sprite[0][34][95] = 1;dino_sprite[0][34][96] = 1;dino_sprite[0][34][97] = 1;dino_sprite[0][34][98] = 1;dino_sprite[0][34][99] = 1;dino_sprite[0][35][44] = 1;dino_sprite[0][35][45] = 1;dino_sprite[0][35][46] = 1;dino_sprite[0][35][47] = 1;dino_sprite[0][35][48] = 1;dino_sprite[0][35][49] = 1;dino_sprite[0][35][50] = 1;dino_sprite[0][35][51] = 1;dino_sprite[0][35][52] = 1;dino_sprite[0][35][53] = 1;dino_sprite[0][35][54] = 1;dino_sprite[0][35][55] = 1;dino_sprite[0][35][56] = 1;dino_sprite[0][35][57] = 1;dino_sprite[0][35][58] = 1;dino_sprite[0][35][59] = 1;dino_sprite[0][35][60] = 1;dino_sprite[0][35][61] = 1;dino_sprite[0][35][62] = 1;dino_sprite[0][35][63] = 1;dino_sprite[0][35][64] = 1;dino_sprite[0][35][65] = 1;dino_sprite[0][35][66] = 1;dino_sprite[0][35][67] = 1;dino_sprite[0][35][68] = 1;dino_sprite[0][35][69] = 1;dino_sprite[0][35][70] = 1;dino_sprite[0][35][71] = 1;dino_sprite[0][35][72] = 1;dino_sprite[0][35][73] = 1;dino_sprite[0][35][74] = 1;dino_sprite[0][35][75] = 1;dino_sprite[0][35][76] = 1;dino_sprite[0][35][77] = 1;dino_sprite[0][35][78] = 1;dino_sprite[0][35][79] = 1;dino_sprite[0][35][80] = 1;dino_sprite[0][35][81] = 1;dino_sprite[0][35][82] = 1;dino_sprite[0][35][83] = 1;dino_sprite[0][35][84] = 1;dino_sprite[0][35][85] = 1;dino_sprite[0][35][86] = 1;dino_sprite[0][35][95] = 1;dino_sprite[0][35][96] = 1;dino_sprite[0][35][97] = 1;dino_sprite[0][35][98] = 1;dino_sprite[0][35][99] = 1;dino_sprite[0][36][44] = 1;dino_sprite[0][36][45] = 1;dino_sprite[0][36][46] = 1;dino_sprite[0][36][47] = 1;dino_sprite[0][36][48] = 1;dino_sprite[0][36][49] = 1;dino_sprite[0][36][50] = 1;dino_sprite[0][36][51] = 1;dino_sprite[0][36][52] = 1;dino_sprite[0][36][53] = 1;dino_sprite[0][36][54] = 1;dino_sprite[0][36][55] = 1;dino_sprite[0][36][56] = 1;dino_sprite[0][36][57] = 1;dino_sprite[0][36][58] = 1;dino_sprite[0][36][59] = 1;dino_sprite[0][36][60] = 1;dino_sprite[0][36][61] = 1;dino_sprite[0][36][62] = 1;dino_sprite[0][36][63] = 1;dino_sprite[0][36][64] = 1;dino_sprite[0][36][65] = 1;dino_sprite[0][36][66] = 1;dino_sprite[0][36][67] = 1;dino_sprite[0][36][68] = 1;dino_sprite[0][36][69] = 1;dino_sprite[0][36][70] = 1;dino_sprite[0][36][71] = 1;dino_sprite[0][36][72] = 1;dino_sprite[0][36][73] = 1;dino_sprite[0][36][74] = 1;dino_sprite[0][36][75] = 1;dino_sprite[0][36][76] = 1;dino_sprite[0][36][77] = 1;dino_sprite[0][36][78] = 1;dino_sprite[0][36][79] = 1;dino_sprite[0][36][80] = 1;dino_sprite[0][36][81] = 1;dino_sprite[0][36][82] = 1;dino_sprite[0][36][83] = 1;dino_sprite[0][36][84] = 1;dino_sprite[0][36][85] = 1;dino_sprite[0][36][86] = 1;dino_sprite[0][36][95] = 1;dino_sprite[0][36][96] = 1;dino_sprite[0][36][97] = 1;dino_sprite[0][36][98] = 1;dino_sprite[0][36][99] = 1;dino_sprite[0][37][44] = 1;dino_sprite[0][37][45] = 1;dino_sprite[0][37][46] = 1;dino_sprite[0][37][47] = 1;dino_sprite[0][37][48] = 1;dino_sprite[0][37][49] = 1;dino_sprite[0][37][50] = 1;dino_sprite[0][37][51] = 1;dino_sprite[0][37][52] = 1;dino_sprite[0][37][53] = 1;dino_sprite[0][37][54] = 1;dino_sprite[0][37][55] = 1;dino_sprite[0][37][56] = 1;dino_sprite[0][37][57] = 1;dino_sprite[0][37][58] = 1;dino_sprite[0][37][59] = 1;dino_sprite[0][37][60] = 1;dino_sprite[0][37][61] = 1;dino_sprite[0][37][62] = 1;dino_sprite[0][37][63] = 1;dino_sprite[0][37][64] = 1;dino_sprite[0][37][65] = 1;dino_sprite[0][37][66] = 1;dino_sprite[0][37][67] = 1;dino_sprite[0][37][68] = 1;dino_sprite[0][37][69] = 1;dino_sprite[0][37][70] = 1;dino_sprite[0][37][71] = 1;dino_sprite[0][37][72] = 1;dino_sprite[0][37][73] = 1;dino_sprite[0][37][74] = 1;dino_sprite[0][37][75] = 1;dino_sprite[0][37][76] = 1;dino_sprite[0][37][77] = 1;dino_sprite[0][37][78] = 1;dino_sprite[0][37][79] = 1;dino_sprite[0][37][80] = 1;dino_sprite[0][37][81] = 1;dino_sprite[0][37][82] = 1;dino_sprite[0][37][83] = 1;dino_sprite[0][37][84] = 1;dino_sprite[0][37][85] = 1;dino_sprite[0][37][86] = 1;dino_sprite[0][38][44] = 1;dino_sprite[0][38][45] = 1;dino_sprite[0][38][46] = 1;dino_sprite[0][38][47] = 1;dino_sprite[0][38][48] = 1;dino_sprite[0][38][49] = 1;dino_sprite[0][38][50] = 1;dino_sprite[0][38][51] = 1;dino_sprite[0][38][52] = 1;dino_sprite[0][38][53] = 1;dino_sprite[0][38][54] = 1;dino_sprite[0][38][55] = 1;dino_sprite[0][38][56] = 1;dino_sprite[0][38][57] = 1;dino_sprite[0][38][58] = 1;dino_sprite[0][38][59] = 1;dino_sprite[0][38][60] = 1;dino_sprite[0][38][61] = 1;dino_sprite[0][38][62] = 1;dino_sprite[0][38][63] = 1;dino_sprite[0][38][64] = 1;dino_sprite[0][38][65] = 1;dino_sprite[0][38][66] = 1;dino_sprite[0][38][67] = 1;dino_sprite[0][38][68] = 1;dino_sprite[0][38][69] = 1;dino_sprite[0][38][70] = 1;dino_sprite[0][38][71] = 1;dino_sprite[0][38][72] = 1;dino_sprite[0][38][73] = 1;dino_sprite[0][38][74] = 1;dino_sprite[0][38][75] = 1;dino_sprite[0][38][76] = 1;dino_sprite[0][38][77] = 1;dino_sprite[0][38][78] = 1;dino_sprite[0][38][79] = 1;dino_sprite[0][38][80] = 1;dino_sprite[0][38][81] = 1;dino_sprite[0][38][82] = 1;dino_sprite[0][38][83] = 1;dino_sprite[0][38][84] = 1;dino_sprite[0][38][85] = 1;dino_sprite[0][38][86] = 1;dino_sprite[0][39][39] = 1;dino_sprite[0][39][40] = 1;dino_sprite[0][39][41] = 1;dino_sprite[0][39][42] = 1;dino_sprite[0][39][43] = 1;dino_sprite[0][39][44] = 1;dino_sprite[0][39][45] = 1;dino_sprite[0][39][46] = 1;dino_sprite[0][39][47] = 1;dino_sprite[0][39][48] = 1;dino_sprite[0][39][49] = 1;dino_sprite[0][39][50] = 1;dino_sprite[0][39][51] = 1;dino_sprite[0][39][52] = 1;dino_sprite[0][39][53] = 1;dino_sprite[0][39][54] = 1;dino_sprite[0][39][55] = 1;dino_sprite[0][39][56] = 1;dino_sprite[0][39][57] = 1;dino_sprite[0][39][58] = 1;dino_sprite[0][39][59] = 1;dino_sprite[0][39][60] = 1;dino_sprite[0][39][61] = 1;dino_sprite[0][39][62] = 1;dino_sprite[0][39][63] = 1;dino_sprite[0][39][64] = 1;dino_sprite[0][39][65] = 1;dino_sprite[0][39][66] = 1;dino_sprite[0][39][67] = 1;dino_sprite[0][39][68] = 1;dino_sprite[0][39][69] = 1;dino_sprite[0][39][70] = 1;dino_sprite[0][39][71] = 1;dino_sprite[0][39][72] = 1;dino_sprite[0][39][73] = 1;dino_sprite[0][39][74] = 1;dino_sprite[0][39][75] = 1;dino_sprite[0][39][76] = 1;dino_sprite[0][39][77] = 1;dino_sprite[0][39][78] = 1;dino_sprite[0][39][79] = 1;dino_sprite[0][39][80] = 1;dino_sprite[0][39][81] = 1;dino_sprite[0][39][82] = 1;dino_sprite[0][39][83] = 1;dino_sprite[0][39][84] = 1;dino_sprite[0][39][85] = 1;dino_sprite[0][39][86] = 1;dino_sprite[0][40][39] = 1;dino_sprite[0][40][40] = 1;dino_sprite[0][40][41] = 1;dino_sprite[0][40][42] = 1;dino_sprite[0][40][43] = 1;dino_sprite[0][40][44] = 1;dino_sprite[0][40][45] = 1;dino_sprite[0][40][46] = 1;dino_sprite[0][40][47] = 1;dino_sprite[0][40][48] = 1;dino_sprite[0][40][49] = 1;dino_sprite[0][40][50] = 1;dino_sprite[0][40][51] = 1;dino_sprite[0][40][52] = 1;dino_sprite[0][40][53] = 1;dino_sprite[0][40][54] = 1;dino_sprite[0][40][55] = 1;dino_sprite[0][40][56] = 1;dino_sprite[0][40][57] = 1;dino_sprite[0][40][58] = 1;dino_sprite[0][40][59] = 1;dino_sprite[0][40][60] = 1;dino_sprite[0][40][61] = 1;dino_sprite[0][40][62] = 1;dino_sprite[0][40][63] = 1;dino_sprite[0][40][64] = 1;dino_sprite[0][40][65] = 1;dino_sprite[0][40][66] = 1;dino_sprite[0][40][67] = 1;dino_sprite[0][40][68] = 1;dino_sprite[0][40][69] = 1;dino_sprite[0][40][70] = 1;dino_sprite[0][40][71] = 1;dino_sprite[0][40][72] = 1;dino_sprite[0][40][73] = 1;dino_sprite[0][40][74] = 1;dino_sprite[0][40][75] = 1;dino_sprite[0][40][76] = 1;dino_sprite[0][40][77] = 1;dino_sprite[0][40][78] = 1;dino_sprite[0][40][79] = 1;dino_sprite[0][40][80] = 1;dino_sprite[0][40][81] = 1;dino_sprite[0][40][82] = 1;dino_sprite[0][40][83] = 1;dino_sprite[0][40][84] = 1;dino_sprite[0][40][85] = 1;dino_sprite[0][40][86] = 1;dino_sprite[0][41][39] = 1;dino_sprite[0][41][40] = 1;dino_sprite[0][41][41] = 1;dino_sprite[0][41][42] = 1;dino_sprite[0][41][43] = 1;dino_sprite[0][41][44] = 1;dino_sprite[0][41][45] = 1;dino_sprite[0][41][46] = 1;dino_sprite[0][41][47] = 1;dino_sprite[0][41][48] = 1;dino_sprite[0][41][49] = 1;dino_sprite[0][41][50] = 1;dino_sprite[0][41][51] = 1;dino_sprite[0][41][52] = 1;dino_sprite[0][41][53] = 1;dino_sprite[0][41][54] = 1;dino_sprite[0][41][55] = 1;dino_sprite[0][41][56] = 1;dino_sprite[0][41][57] = 1;dino_sprite[0][41][58] = 1;dino_sprite[0][41][59] = 1;dino_sprite[0][41][60] = 1;dino_sprite[0][41][61] = 1;dino_sprite[0][41][62] = 1;dino_sprite[0][41][63] = 1;dino_sprite[0][41][64] = 1;dino_sprite[0][41][65] = 1;dino_sprite[0][41][66] = 1;dino_sprite[0][41][67] = 1;dino_sprite[0][41][68] = 1;dino_sprite[0][41][69] = 1;dino_sprite[0][41][70] = 1;dino_sprite[0][41][71] = 1;dino_sprite[0][41][72] = 1;dino_sprite[0][41][73] = 1;dino_sprite[0][41][74] = 1;dino_sprite[0][41][75] = 1;dino_sprite[0][41][76] = 1;dino_sprite[0][41][77] = 1;dino_sprite[0][41][78] = 1;dino_sprite[0][41][79] = 1;dino_sprite[0][41][80] = 1;dino_sprite[0][41][81] = 1;dino_sprite[0][41][82] = 1;dino_sprite[0][42][39] = 1;dino_sprite[0][42][40] = 1;dino_sprite[0][42][41] = 1;dino_sprite[0][42][42] = 1;dino_sprite[0][42][43] = 1;dino_sprite[0][42][44] = 1;dino_sprite[0][42][45] = 1;dino_sprite[0][42][46] = 1;dino_sprite[0][42][47] = 1;dino_sprite[0][42][48] = 1;dino_sprite[0][42][49] = 1;dino_sprite[0][42][50] = 1;dino_sprite[0][42][51] = 1;dino_sprite[0][42][52] = 1;dino_sprite[0][42][53] = 1;dino_sprite[0][42][54] = 1;dino_sprite[0][42][55] = 1;dino_sprite[0][42][56] = 1;dino_sprite[0][42][57] = 1;dino_sprite[0][42][58] = 1;dino_sprite[0][42][59] = 1;dino_sprite[0][42][60] = 1;dino_sprite[0][42][61] = 1;dino_sprite[0][42][62] = 1;dino_sprite[0][42][63] = 1;dino_sprite[0][42][64] = 1;dino_sprite[0][42][65] = 1;dino_sprite[0][42][66] = 1;dino_sprite[0][42][67] = 1;dino_sprite[0][42][68] = 1;dino_sprite[0][42][69] = 1;dino_sprite[0][42][70] = 1;dino_sprite[0][42][71] = 1;dino_sprite[0][42][72] = 1;dino_sprite[0][42][73] = 1;dino_sprite[0][42][74] = 1;dino_sprite[0][42][75] = 1;dino_sprite[0][42][76] = 1;dino_sprite[0][42][77] = 1;dino_sprite[0][42][78] = 1;dino_sprite[0][42][79] = 1;dino_sprite[0][42][80] = 1;dino_sprite[0][42][81] = 1;dino_sprite[0][42][82] = 1;dino_sprite[0][43][39] = 1;dino_sprite[0][43][40] = 1;dino_sprite[0][43][41] = 1;dino_sprite[0][43][42] = 1;dino_sprite[0][43][43] = 1;dino_sprite[0][43][44] = 1;dino_sprite[0][43][45] = 1;dino_sprite[0][43][46] = 1;dino_sprite[0][43][47] = 1;dino_sprite[0][43][48] = 1;dino_sprite[0][43][49] = 1;dino_sprite[0][43][50] = 1;dino_sprite[0][43][51] = 1;dino_sprite[0][43][52] = 1;dino_sprite[0][43][53] = 1;dino_sprite[0][43][54] = 1;dino_sprite[0][43][55] = 1;dino_sprite[0][43][56] = 1;dino_sprite[0][43][57] = 1;dino_sprite[0][43][58] = 1;dino_sprite[0][43][59] = 1;dino_sprite[0][43][60] = 1;dino_sprite[0][43][61] = 1;dino_sprite[0][43][62] = 1;dino_sprite[0][43][63] = 1;dino_sprite[0][43][64] = 1;dino_sprite[0][43][65] = 1;dino_sprite[0][43][66] = 1;dino_sprite[0][43][67] = 1;dino_sprite[0][43][68] = 1;dino_sprite[0][43][69] = 1;dino_sprite[0][43][70] = 1;dino_sprite[0][43][71] = 1;dino_sprite[0][43][72] = 1;dino_sprite[0][43][73] = 1;dino_sprite[0][43][74] = 1;dino_sprite[0][43][75] = 1;dino_sprite[0][43][76] = 1;dino_sprite[0][43][77] = 1;dino_sprite[0][43][78] = 1;dino_sprite[0][43][79] = 1;dino_sprite[0][43][80] = 1;dino_sprite[0][43][81] = 1;dino_sprite[0][43][82] = 1;dino_sprite[0][44][39] = 1;dino_sprite[0][44][40] = 1;dino_sprite[0][44][41] = 1;dino_sprite[0][44][42] = 1;dino_sprite[0][44][43] = 1;dino_sprite[0][44][44] = 1;dino_sprite[0][44][45] = 1;dino_sprite[0][44][46] = 1;dino_sprite[0][44][47] = 1;dino_sprite[0][44][48] = 1;dino_sprite[0][44][49] = 1;dino_sprite[0][44][50] = 1;dino_sprite[0][44][51] = 1;dino_sprite[0][44][52] = 1;dino_sprite[0][44][53] = 1;dino_sprite[0][44][54] = 1;dino_sprite[0][44][55] = 1;dino_sprite[0][44][56] = 1;dino_sprite[0][44][57] = 1;dino_sprite[0][44][58] = 1;dino_sprite[0][44][59] = 1;dino_sprite[0][44][60] = 1;dino_sprite[0][44][61] = 1;dino_sprite[0][44][62] = 1;dino_sprite[0][44][63] = 1;dino_sprite[0][44][64] = 1;dino_sprite[0][44][65] = 1;dino_sprite[0][44][66] = 1;dino_sprite[0][44][67] = 1;dino_sprite[0][44][68] = 1;dino_sprite[0][44][69] = 1;dino_sprite[0][44][70] = 1;dino_sprite[0][44][71] = 1;dino_sprite[0][44][72] = 1;dino_sprite[0][44][73] = 1;dino_sprite[0][44][74] = 1;dino_sprite[0][44][75] = 1;dino_sprite[0][44][76] = 1;dino_sprite[0][44][77] = 1;dino_sprite[0][44][78] = 1;dino_sprite[0][44][79] = 1;dino_sprite[0][44][80] = 1;dino_sprite[0][44][81] = 1;dino_sprite[0][44][82] = 1;dino_sprite[0][45][35] = 1;dino_sprite[0][45][36] = 1;dino_sprite[0][45][37] = 1;dino_sprite[0][45][39] = 1;dino_sprite[0][45][40] = 1;dino_sprite[0][45][41] = 1;dino_sprite[0][45][42] = 1;dino_sprite[0][45][43] = 1;dino_sprite[0][45][44] = 1;dino_sprite[0][45][45] = 1;dino_sprite[0][45][46] = 1;dino_sprite[0][45][47] = 1;dino_sprite[0][45][48] = 1;dino_sprite[0][45][49] = 1;dino_sprite[0][45][50] = 1;dino_sprite[0][45][51] = 1;dino_sprite[0][45][52] = 1;dino_sprite[0][45][53] = 1;dino_sprite[0][45][54] = 1;dino_sprite[0][45][55] = 1;dino_sprite[0][45][56] = 1;dino_sprite[0][45][57] = 1;dino_sprite[0][45][58] = 1;dino_sprite[0][45][59] = 1;dino_sprite[0][45][60] = 1;dino_sprite[0][45][61] = 1;dino_sprite[0][45][62] = 1;dino_sprite[0][45][63] = 1;dino_sprite[0][45][64] = 1;dino_sprite[0][45][65] = 1;dino_sprite[0][45][66] = 1;dino_sprite[0][45][67] = 1;dino_sprite[0][45][68] = 1;dino_sprite[0][45][69] = 1;dino_sprite[0][45][70] = 1;dino_sprite[0][45][71] = 1;dino_sprite[0][45][72] = 1;dino_sprite[0][45][73] = 1;dino_sprite[0][45][74] = 1;dino_sprite[0][45][75] = 1;dino_sprite[0][45][76] = 1;dino_sprite[0][45][77] = 1;dino_sprite[0][45][78] = 1;dino_sprite[0][45][79] = 1;dino_sprite[0][45][80] = 1;dino_sprite[0][45][81] = 1;dino_sprite[0][45][82] = 1;dino_sprite[0][45][84] = 1;dino_sprite[0][45][85] = 1;dino_sprite[0][45][86] = 1;dino_sprite[0][46][35] = 1;dino_sprite[0][46][36] = 1;dino_sprite[0][46][37] = 1;dino_sprite[0][46][38] = 1;dino_sprite[0][46][39] = 1;dino_sprite[0][46][40] = 1;dino_sprite[0][46][41] = 1;dino_sprite[0][46][42] = 1;dino_sprite[0][46][43] = 1;dino_sprite[0][46][44] = 1;dino_sprite[0][46][45] = 1;dino_sprite[0][46][46] = 1;dino_sprite[0][46][47] = 1;dino_sprite[0][46][48] = 1;dino_sprite[0][46][49] = 1;dino_sprite[0][46][50] = 1;dino_sprite[0][46][51] = 1;dino_sprite[0][46][52] = 1;dino_sprite[0][46][53] = 1;dino_sprite[0][46][54] = 1;dino_sprite[0][46][55] = 1;dino_sprite[0][46][56] = 1;dino_sprite[0][46][57] = 1;dino_sprite[0][46][58] = 1;dino_sprite[0][46][59] = 1;dino_sprite[0][46][60] = 1;dino_sprite[0][46][61] = 1;dino_sprite[0][46][62] = 1;dino_sprite[0][46][63] = 1;dino_sprite[0][46][64] = 1;dino_sprite[0][46][65] = 1;dino_sprite[0][46][66] = 1;dino_sprite[0][46][67] = 1;dino_sprite[0][46][68] = 1;dino_sprite[0][46][69] = 1;dino_sprite[0][46][70] = 1;dino_sprite[0][46][71] = 1;dino_sprite[0][46][72] = 1;dino_sprite[0][46][73] = 1;dino_sprite[0][46][74] = 1;dino_sprite[0][46][75] = 1;dino_sprite[0][46][76] = 1;dino_sprite[0][46][77] = 1;dino_sprite[0][46][78] = 1;dino_sprite[0][46][79] = 1;dino_sprite[0][46][80] = 1;dino_sprite[0][46][81] = 1;dino_sprite[0][46][82] = 1;dino_sprite[0][46][83] = 1;dino_sprite[0][46][84] = 1;dino_sprite[0][46][85] = 1;dino_sprite[0][46][86] = 1;dino_sprite[0][47][35] = 1;dino_sprite[0][47][36] = 1;dino_sprite[0][47][37] = 1;dino_sprite[0][47][38] = 1;dino_sprite[0][47][39] = 1;dino_sprite[0][47][40] = 1;dino_sprite[0][47][41] = 1;dino_sprite[0][47][42] = 1;dino_sprite[0][47][43] = 1;dino_sprite[0][47][44] = 1;dino_sprite[0][47][45] = 1;dino_sprite[0][47][46] = 1;dino_sprite[0][47][47] = 1;dino_sprite[0][47][48] = 1;dino_sprite[0][47][49] = 1;dino_sprite[0][47][50] = 1;dino_sprite[0][47][51] = 1;dino_sprite[0][47][52] = 1;dino_sprite[0][47][53] = 1;dino_sprite[0][47][54] = 1;dino_sprite[0][47][55] = 1;dino_sprite[0][47][56] = 1;dino_sprite[0][47][57] = 1;dino_sprite[0][47][58] = 1;dino_sprite[0][47][59] = 1;dino_sprite[0][47][60] = 1;dino_sprite[0][47][61] = 1;dino_sprite[0][47][62] = 1;dino_sprite[0][47][63] = 1;dino_sprite[0][47][64] = 1;dino_sprite[0][47][65] = 1;dino_sprite[0][47][66] = 1;dino_sprite[0][47][67] = 1;dino_sprite[0][47][68] = 1;dino_sprite[0][47][69] = 1;dino_sprite[0][47][70] = 1;dino_sprite[0][47][71] = 1;dino_sprite[0][47][72] = 1;dino_sprite[0][47][73] = 1;dino_sprite[0][47][74] = 1;dino_sprite[0][47][75] = 1;dino_sprite[0][47][76] = 1;dino_sprite[0][47][77] = 1;dino_sprite[0][47][78] = 1;dino_sprite[0][47][79] = 1;dino_sprite[0][47][80] = 1;dino_sprite[0][47][81] = 1;dino_sprite[0][47][82] = 1;dino_sprite[0][47][83] = 1;dino_sprite[0][47][84] = 1;dino_sprite[0][47][85] = 1;dino_sprite[0][47][86] = 1;dino_sprite[0][48][35] = 1;dino_sprite[0][48][36] = 1;dino_sprite[0][48][37] = 1;dino_sprite[0][48][38] = 1;dino_sprite[0][48][39] = 1;dino_sprite[0][48][40] = 1;dino_sprite[0][48][41] = 1;dino_sprite[0][48][42] = 1;dino_sprite[0][48][43] = 1;dino_sprite[0][48][44] = 1;dino_sprite[0][48][45] = 1;dino_sprite[0][48][46] = 1;dino_sprite[0][48][47] = 1;dino_sprite[0][48][48] = 1;dino_sprite[0][48][49] = 1;dino_sprite[0][48][50] = 1;dino_sprite[0][48][51] = 1;dino_sprite[0][48][52] = 1;dino_sprite[0][48][53] = 1;dino_sprite[0][48][54] = 1;dino_sprite[0][48][55] = 1;dino_sprite[0][48][56] = 1;dino_sprite[0][48][57] = 1;dino_sprite[0][48][58] = 1;dino_sprite[0][48][59] = 1;dino_sprite[0][48][60] = 1;dino_sprite[0][48][61] = 1;dino_sprite[0][48][62] = 1;dino_sprite[0][48][63] = 1;dino_sprite[0][48][64] = 1;dino_sprite[0][48][65] = 1;dino_sprite[0][48][66] = 1;dino_sprite[0][48][67] = 1;dino_sprite[0][48][68] = 1;dino_sprite[0][48][69] = 1;dino_sprite[0][48][70] = 1;dino_sprite[0][48][71] = 1;dino_sprite[0][48][72] = 1;dino_sprite[0][48][73] = 1;dino_sprite[0][48][74] = 1;dino_sprite[0][48][75] = 1;dino_sprite[0][48][76] = 1;dino_sprite[0][48][77] = 1;dino_sprite[0][48][78] = 1;dino_sprite[0][48][79] = 1;dino_sprite[0][48][80] = 1;dino_sprite[0][48][81] = 1;dino_sprite[0][48][82] = 1;dino_sprite[0][48][83] = 1;dino_sprite[0][48][84] = 1;dino_sprite[0][48][85] = 1;dino_sprite[0][48][86] = 1;dino_sprite[0][49][35] = 1;dino_sprite[0][49][36] = 1;dino_sprite[0][49][37] = 1;dino_sprite[0][49][38] = 1;dino_sprite[0][49][39] = 1;dino_sprite[0][49][40] = 1;dino_sprite[0][49][41] = 1;dino_sprite[0][49][42] = 1;dino_sprite[0][49][43] = 1;dino_sprite[0][49][44] = 1;dino_sprite[0][49][45] = 1;dino_sprite[0][49][46] = 1;dino_sprite[0][49][47] = 1;dino_sprite[0][49][48] = 1;dino_sprite[0][49][49] = 1;dino_sprite[0][49][50] = 1;dino_sprite[0][49][51] = 1;dino_sprite[0][49][52] = 1;dino_sprite[0][49][53] = 1;dino_sprite[0][49][54] = 1;dino_sprite[0][49][55] = 1;dino_sprite[0][49][56] = 1;dino_sprite[0][49][57] = 1;dino_sprite[0][49][58] = 1;dino_sprite[0][49][59] = 1;dino_sprite[0][49][60] = 1;dino_sprite[0][49][61] = 1;dino_sprite[0][49][62] = 1;dino_sprite[0][49][63] = 1;dino_sprite[0][49][64] = 1;dino_sprite[0][49][65] = 1;dino_sprite[0][49][66] = 1;dino_sprite[0][49][67] = 1;dino_sprite[0][49][68] = 1;dino_sprite[0][49][69] = 1;dino_sprite[0][49][70] = 1;dino_sprite[0][49][71] = 1;dino_sprite[0][49][72] = 1;dino_sprite[0][49][73] = 1;dino_sprite[0][49][74] = 1;dino_sprite[0][49][75] = 1;dino_sprite[0][49][76] = 1;dino_sprite[0][49][77] = 1;dino_sprite[0][49][78] = 1;dino_sprite[0][49][79] = 1;dino_sprite[0][49][80] = 1;dino_sprite[0][49][81] = 1;dino_sprite[0][49][82] = 1;dino_sprite[0][49][83] = 1;dino_sprite[0][49][84] = 1;dino_sprite[0][49][85] = 1;dino_sprite[0][49][86] = 1;dino_sprite[0][50][35] = 1;dino_sprite[0][50][36] = 1;dino_sprite[0][50][37] = 1;dino_sprite[0][50][38] = 1;dino_sprite[0][50][39] = 1;dino_sprite[0][50][40] = 1;dino_sprite[0][50][41] = 1;dino_sprite[0][50][42] = 1;dino_sprite[0][50][43] = 1;dino_sprite[0][50][44] = 1;dino_sprite[0][50][45] = 1;dino_sprite[0][50][46] = 1;dino_sprite[0][50][47] = 1;dino_sprite[0][50][48] = 1;dino_sprite[0][50][49] = 1;dino_sprite[0][50][50] = 1;dino_sprite[0][50][51] = 1;dino_sprite[0][50][52] = 1;dino_sprite[0][50][53] = 1;dino_sprite[0][50][54] = 1;dino_sprite[0][50][55] = 1;dino_sprite[0][50][56] = 1;dino_sprite[0][50][57] = 1;dino_sprite[0][50][58] = 1;dino_sprite[0][50][59] = 1;dino_sprite[0][50][60] = 1;dino_sprite[0][50][61] = 1;dino_sprite[0][50][62] = 1;dino_sprite[0][50][63] = 1;dino_sprite[0][50][64] = 1;dino_sprite[0][50][65] = 1;dino_sprite[0][50][66] = 1;dino_sprite[0][50][67] = 1;dino_sprite[0][50][68] = 1;dino_sprite[0][50][69] = 1;dino_sprite[0][50][70] = 1;dino_sprite[0][50][71] = 1;dino_sprite[0][50][72] = 1;dino_sprite[0][50][73] = 1;dino_sprite[0][50][74] = 1;dino_sprite[0][50][75] = 1;dino_sprite[0][50][76] = 1;dino_sprite[0][50][77] = 1;dino_sprite[0][50][78] = 1;dino_sprite[0][50][79] = 1;dino_sprite[0][50][80] = 1;dino_sprite[0][50][81] = 1;dino_sprite[0][50][82] = 1;dino_sprite[0][50][83] = 1;dino_sprite[0][50][84] = 1;dino_sprite[0][50][85] = 1;dino_sprite[0][50][86] = 1;dino_sprite[0][50][88] = 1;dino_sprite[0][50][89] = 1;dino_sprite[0][50][90] = 1;dino_sprite[0][50][91] = 1;dino_sprite[0][50][92] = 1;dino_sprite[0][50][93] = 1;dino_sprite[0][50][94] = 1;dino_sprite[0][50][95] = 1;dino_sprite[0][50][96] = 1;dino_sprite[0][50][97] = 1;dino_sprite[0][50][98] = 1;dino_sprite[0][50][99] = 1;dino_sprite[0][51][3] = 1;dino_sprite[0][51][4] = 1;dino_sprite[0][51][5] = 1;dino_sprite[0][51][6] = 1;dino_sprite[0][51][7] = 1;dino_sprite[0][51][8] = 1;dino_sprite[0][51][9] = 1;dino_sprite[0][51][10] = 1;dino_sprite[0][51][11] = 1;dino_sprite[0][51][12] = 1;dino_sprite[0][51][13] = 1;dino_sprite[0][51][14] = 1;dino_sprite[0][51][15] = 1;dino_sprite[0][51][16] = 1;dino_sprite[0][51][17] = 1;dino_sprite[0][51][18] = 1;dino_sprite[0][51][19] = 1;dino_sprite[0][51][20] = 1;dino_sprite[0][51][21] = 1;dino_sprite[0][51][22] = 1;dino_sprite[0][51][23] = 1;dino_sprite[0][51][24] = 1;dino_sprite[0][51][25] = 1;dino_sprite[0][51][26] = 1;dino_sprite[0][51][27] = 1;dino_sprite[0][51][28] = 1;dino_sprite[0][51][29] = 1;dino_sprite[0][51][30] = 1;dino_sprite[0][51][31] = 1;dino_sprite[0][51][32] = 1;dino_sprite[0][51][33] = 1;dino_sprite[0][51][34] = 1;dino_sprite[0][51][35] = 1;dino_sprite[0][51][36] = 1;dino_sprite[0][51][37] = 1;dino_sprite[0][51][38] = 1;dino_sprite[0][51][39] = 1;dino_sprite[0][51][40] = 1;dino_sprite[0][51][41] = 1;dino_sprite[0][51][42] = 1;dino_sprite[0][51][43] = 1;dino_sprite[0][51][44] = 1;dino_sprite[0][51][45] = 1;dino_sprite[0][51][46] = 1;dino_sprite[0][51][47] = 1;dino_sprite[0][51][48] = 1;dino_sprite[0][51][49] = 1;dino_sprite[0][51][50] = 1;dino_sprite[0][51][51] = 1;dino_sprite[0][51][52] = 1;dino_sprite[0][51][53] = 1;dino_sprite[0][51][54] = 1;dino_sprite[0][51][55] = 1;dino_sprite[0][51][56] = 1;dino_sprite[0][51][57] = 1;dino_sprite[0][51][58] = 1;dino_sprite[0][51][59] = 1;dino_sprite[0][51][60] = 1;dino_sprite[0][51][61] = 1;dino_sprite[0][51][62] = 1;dino_sprite[0][51][63] = 1;dino_sprite[0][51][64] = 1;dino_sprite[0][51][65] = 1;dino_sprite[0][51][66] = 1;dino_sprite[0][51][67] = 1;dino_sprite[0][51][68] = 1;dino_sprite[0][51][69] = 1;dino_sprite[0][51][70] = 1;dino_sprite[0][51][71] = 1;dino_sprite[0][51][72] = 1;dino_sprite[0][51][73] = 1;dino_sprite[0][51][74] = 1;dino_sprite[0][51][75] = 1;dino_sprite[0][51][76] = 1;dino_sprite[0][51][77] = 1;dino_sprite[0][51][78] = 1;dino_sprite[0][51][79] = 1;dino_sprite[0][51][80] = 1;dino_sprite[0][51][81] = 1;dino_sprite[0][51][82] = 1;dino_sprite[0][51][83] = 1;dino_sprite[0][51][84] = 1;dino_sprite[0][51][85] = 1;dino_sprite[0][51][86] = 1;dino_sprite[0][51][87] = 1;dino_sprite[0][51][88] = 1;dino_sprite[0][51][89] = 1;dino_sprite[0][51][90] = 1;dino_sprite[0][51][91] = 1;dino_sprite[0][51][92] = 1;dino_sprite[0][51][93] = 1;dino_sprite[0][51][94] = 1;dino_sprite[0][51][95] = 1;dino_sprite[0][51][96] = 1;dino_sprite[0][51][97] = 1;dino_sprite[0][51][98] = 1;dino_sprite[0][51][99] = 1;dino_sprite[0][52][3] = 1;dino_sprite[0][52][4] = 1;dino_sprite[0][52][5] = 1;dino_sprite[0][52][6] = 1;dino_sprite[0][52][7] = 1;dino_sprite[0][52][8] = 1;dino_sprite[0][52][9] = 1;dino_sprite[0][52][10] = 1;dino_sprite[0][52][11] = 1;dino_sprite[0][52][12] = 1;dino_sprite[0][52][13] = 1;dino_sprite[0][52][14] = 1;dino_sprite[0][52][15] = 1;dino_sprite[0][52][16] = 1;dino_sprite[0][52][17] = 1;dino_sprite[0][52][18] = 1;dino_sprite[0][52][19] = 1;dino_sprite[0][52][20] = 1;dino_sprite[0][52][21] = 1;dino_sprite[0][52][22] = 1;dino_sprite[0][52][23] = 1;dino_sprite[0][52][24] = 1;dino_sprite[0][52][25] = 1;dino_sprite[0][52][26] = 1;dino_sprite[0][52][27] = 1;dino_sprite[0][52][28] = 1;dino_sprite[0][52][29] = 1;dino_sprite[0][52][30] = 1;dino_sprite[0][52][31] = 1;dino_sprite[0][52][32] = 1;dino_sprite[0][52][33] = 1;dino_sprite[0][52][34] = 1;dino_sprite[0][52][35] = 1;dino_sprite[0][52][36] = 1;dino_sprite[0][52][37] = 1;dino_sprite[0][52][38] = 1;dino_sprite[0][52][39] = 1;dino_sprite[0][52][40] = 1;dino_sprite[0][52][41] = 1;dino_sprite[0][52][42] = 1;dino_sprite[0][52][43] = 1;dino_sprite[0][52][44] = 1;dino_sprite[0][52][45] = 1;dino_sprite[0][52][46] = 1;dino_sprite[0][52][47] = 1;dino_sprite[0][52][48] = 1;dino_sprite[0][52][49] = 1;dino_sprite[0][52][50] = 1;dino_sprite[0][52][51] = 1;dino_sprite[0][52][52] = 1;dino_sprite[0][52][53] = 1;dino_sprite[0][52][54] = 1;dino_sprite[0][52][55] = 1;dino_sprite[0][52][56] = 1;dino_sprite[0][52][57] = 1;dino_sprite[0][52][58] = 1;dino_sprite[0][52][59] = 1;dino_sprite[0][52][60] = 1;dino_sprite[0][52][61] = 1;dino_sprite[0][52][62] = 1;dino_sprite[0][52][63] = 1;dino_sprite[0][52][64] = 1;dino_sprite[0][52][65] = 1;dino_sprite[0][52][66] = 1;dino_sprite[0][52][67] = 1;dino_sprite[0][52][68] = 1;dino_sprite[0][52][69] = 1;dino_sprite[0][52][70] = 1;dino_sprite[0][52][71] = 1;dino_sprite[0][52][72] = 1;dino_sprite[0][52][73] = 1;dino_sprite[0][52][74] = 1;dino_sprite[0][52][75] = 1;dino_sprite[0][52][76] = 1;dino_sprite[0][52][77] = 1;dino_sprite[0][52][78] = 1;dino_sprite[0][52][79] = 1;dino_sprite[0][52][80] = 1;dino_sprite[0][52][81] = 1;dino_sprite[0][52][82] = 1;dino_sprite[0][52][83] = 1;dino_sprite[0][52][84] = 1;dino_sprite[0][52][85] = 1;dino_sprite[0][52][86] = 1;dino_sprite[0][52][87] = 1;dino_sprite[0][52][88] = 1;dino_sprite[0][52][89] = 1;dino_sprite[0][52][90] = 1;dino_sprite[0][52][91] = 1;dino_sprite[0][52][92] = 1;dino_sprite[0][52][93] = 1;dino_sprite[0][52][94] = 1;dino_sprite[0][52][95] = 1;dino_sprite[0][52][96] = 1;dino_sprite[0][52][97] = 1;dino_sprite[0][52][98] = 1;dino_sprite[0][52][99] = 1;dino_sprite[0][53][3] = 1;dino_sprite[0][53][4] = 1;dino_sprite[0][53][5] = 1;dino_sprite[0][53][6] = 1;dino_sprite[0][53][7] = 1;dino_sprite[0][53][8] = 1;dino_sprite[0][53][9] = 1;dino_sprite[0][53][10] = 1;dino_sprite[0][53][11] = 1;dino_sprite[0][53][12] = 1;dino_sprite[0][53][13] = 1;dino_sprite[0][53][14] = 1;dino_sprite[0][53][15] = 1;dino_sprite[0][53][16] = 1;dino_sprite[0][53][17] = 1;dino_sprite[0][53][18] = 1;dino_sprite[0][53][19] = 1;dino_sprite[0][53][20] = 1;dino_sprite[0][53][21] = 1;dino_sprite[0][53][22] = 1;dino_sprite[0][53][23] = 1;dino_sprite[0][53][24] = 1;dino_sprite[0][53][25] = 1;dino_sprite[0][53][26] = 1;dino_sprite[0][53][27] = 1;dino_sprite[0][53][28] = 1;dino_sprite[0][53][29] = 1;dino_sprite[0][53][30] = 1;dino_sprite[0][53][31] = 1;dino_sprite[0][53][32] = 1;dino_sprite[0][53][33] = 1;dino_sprite[0][53][34] = 1;dino_sprite[0][53][35] = 1;dino_sprite[0][53][36] = 1;dino_sprite[0][53][37] = 1;dino_sprite[0][53][38] = 1;dino_sprite[0][53][39] = 1;dino_sprite[0][53][40] = 1;dino_sprite[0][53][41] = 1;dino_sprite[0][53][42] = 1;dino_sprite[0][53][43] = 1;dino_sprite[0][53][44] = 1;dino_sprite[0][53][45] = 1;dino_sprite[0][53][46] = 1;dino_sprite[0][53][47] = 1;dino_sprite[0][53][48] = 1;dino_sprite[0][53][49] = 1;dino_sprite[0][53][50] = 1;dino_sprite[0][53][51] = 1;dino_sprite[0][53][52] = 1;dino_sprite[0][53][53] = 1;dino_sprite[0][53][54] = 1;dino_sprite[0][53][55] = 1;dino_sprite[0][53][56] = 1;dino_sprite[0][53][57] = 1;dino_sprite[0][53][58] = 1;dino_sprite[0][53][59] = 1;dino_sprite[0][53][60] = 1;dino_sprite[0][53][61] = 1;dino_sprite[0][53][62] = 1;dino_sprite[0][53][63] = 1;dino_sprite[0][53][64] = 1;dino_sprite[0][53][65] = 1;dino_sprite[0][53][66] = 1;dino_sprite[0][53][67] = 1;dino_sprite[0][53][68] = 1;dino_sprite[0][53][69] = 1;dino_sprite[0][53][70] = 1;dino_sprite[0][53][71] = 1;dino_sprite[0][53][72] = 1;dino_sprite[0][53][73] = 1;dino_sprite[0][53][74] = 1;dino_sprite[0][53][75] = 1;dino_sprite[0][53][76] = 1;dino_sprite[0][53][77] = 1;dino_sprite[0][53][78] = 1;dino_sprite[0][53][79] = 1;dino_sprite[0][53][80] = 1;dino_sprite[0][53][81] = 1;dino_sprite[0][53][82] = 1;dino_sprite[0][53][83] = 1;dino_sprite[0][53][84] = 1;dino_sprite[0][53][85] = 1;dino_sprite[0][53][86] = 1;dino_sprite[0][53][87] = 1;dino_sprite[0][53][88] = 1;dino_sprite[0][53][89] = 1;dino_sprite[0][53][90] = 1;dino_sprite[0][53][91] = 1;dino_sprite[0][53][92] = 1;dino_sprite[0][53][93] = 1;dino_sprite[0][53][94] = 1;dino_sprite[0][53][95] = 1;dino_sprite[0][53][96] = 1;dino_sprite[0][53][97] = 1;dino_sprite[0][53][98] = 1;dino_sprite[0][53][99] = 1;dino_sprite[0][54][3] = 1;dino_sprite[0][54][4] = 1;dino_sprite[0][54][5] = 1;dino_sprite[0][54][6] = 1;dino_sprite[0][54][7] = 1;dino_sprite[0][54][8] = 1;dino_sprite[0][54][9] = 1;dino_sprite[0][54][10] = 1;dino_sprite[0][54][11] = 1;dino_sprite[0][54][12] = 1;dino_sprite[0][54][13] = 1;dino_sprite[0][54][14] = 1;dino_sprite[0][54][15] = 1;dino_sprite[0][54][16] = 1;dino_sprite[0][54][17] = 1;dino_sprite[0][54][18] = 1;dino_sprite[0][54][19] = 1;dino_sprite[0][54][20] = 1;dino_sprite[0][54][21] = 1;dino_sprite[0][54][22] = 1;dino_sprite[0][54][23] = 1;dino_sprite[0][54][24] = 1;dino_sprite[0][54][25] = 1;dino_sprite[0][54][26] = 1;dino_sprite[0][54][27] = 1;dino_sprite[0][54][28] = 1;dino_sprite[0][54][29] = 1;dino_sprite[0][54][30] = 1;dino_sprite[0][54][31] = 1;dino_sprite[0][54][32] = 1;dino_sprite[0][54][33] = 1;dino_sprite[0][54][34] = 1;dino_sprite[0][54][35] = 1;dino_sprite[0][54][36] = 1;dino_sprite[0][54][37] = 1;dino_sprite[0][54][38] = 1;dino_sprite[0][54][39] = 1;dino_sprite[0][54][40] = 1;dino_sprite[0][54][41] = 1;dino_sprite[0][54][42] = 1;dino_sprite[0][54][43] = 1;dino_sprite[0][54][44] = 1;dino_sprite[0][54][45] = 1;dino_sprite[0][54][46] = 1;dino_sprite[0][54][47] = 1;dino_sprite[0][54][48] = 1;dino_sprite[0][54][49] = 1;dino_sprite[0][54][50] = 1;dino_sprite[0][54][51] = 1;dino_sprite[0][54][52] = 1;dino_sprite[0][54][53] = 1;dino_sprite[0][54][54] = 1;dino_sprite[0][54][55] = 1;dino_sprite[0][54][56] = 1;dino_sprite[0][54][57] = 1;dino_sprite[0][54][58] = 1;dino_sprite[0][54][59] = 1;dino_sprite[0][54][60] = 1;dino_sprite[0][54][61] = 1;dino_sprite[0][54][62] = 1;dino_sprite[0][54][63] = 1;dino_sprite[0][54][64] = 1;dino_sprite[0][54][65] = 1;dino_sprite[0][54][66] = 1;dino_sprite[0][54][67] = 1;dino_sprite[0][54][68] = 1;dino_sprite[0][54][69] = 1;dino_sprite[0][54][70] = 1;dino_sprite[0][54][71] = 1;dino_sprite[0][54][72] = 1;dino_sprite[0][54][73] = 1;dino_sprite[0][54][74] = 1;dino_sprite[0][54][75] = 1;dino_sprite[0][54][76] = 1;dino_sprite[0][54][77] = 1;dino_sprite[0][54][78] = 1;dino_sprite[0][54][79] = 1;dino_sprite[0][54][80] = 1;dino_sprite[0][54][81] = 1;dino_sprite[0][54][82] = 1;dino_sprite[0][54][83] = 1;dino_sprite[0][54][84] = 1;dino_sprite[0][54][85] = 1;dino_sprite[0][54][86] = 1;dino_sprite[0][54][87] = 1;dino_sprite[0][54][88] = 1;dino_sprite[0][54][89] = 1;dino_sprite[0][54][90] = 1;dino_sprite[0][54][91] = 1;dino_sprite[0][54][92] = 1;dino_sprite[0][54][93] = 1;dino_sprite[0][54][94] = 1;dino_sprite[0][54][95] = 1;dino_sprite[0][54][96] = 1;dino_sprite[0][54][97] = 1;dino_sprite[0][54][98] = 1;dino_sprite[0][54][99] = 1;dino_sprite[0][55][3] = 1;dino_sprite[0][55][4] = 1;dino_sprite[0][55][5] = 1;dino_sprite[0][55][6] = 1;dino_sprite[0][55][7] = 1;dino_sprite[0][55][8] = 1;dino_sprite[0][55][9] = 1;dino_sprite[0][55][10] = 1;dino_sprite[0][55][11] = 1;dino_sprite[0][55][12] = 1;dino_sprite[0][55][13] = 1;dino_sprite[0][55][14] = 1;dino_sprite[0][55][15] = 1;dino_sprite[0][55][16] = 1;dino_sprite[0][55][17] = 1;dino_sprite[0][55][18] = 1;dino_sprite[0][55][19] = 1;dino_sprite[0][55][20] = 1;dino_sprite[0][55][21] = 1;dino_sprite[0][55][22] = 1;dino_sprite[0][55][23] = 1;dino_sprite[0][55][24] = 1;dino_sprite[0][55][25] = 1;dino_sprite[0][55][26] = 1;dino_sprite[0][55][27] = 1;dino_sprite[0][55][28] = 1;dino_sprite[0][55][29] = 1;dino_sprite[0][55][30] = 1;dino_sprite[0][55][31] = 1;dino_sprite[0][55][32] = 1;dino_sprite[0][55][33] = 1;dino_sprite[0][55][34] = 1;dino_sprite[0][55][35] = 1;dino_sprite[0][55][36] = 1;dino_sprite[0][55][37] = 1;dino_sprite[0][55][38] = 1;dino_sprite[0][55][39] = 1;dino_sprite[0][55][40] = 1;dino_sprite[0][55][41] = 1;dino_sprite[0][55][42] = 1;dino_sprite[0][55][43] = 1;dino_sprite[0][55][44] = 1;dino_sprite[0][55][45] = 1;dino_sprite[0][55][46] = 1;dino_sprite[0][55][47] = 1;dino_sprite[0][55][48] = 1;dino_sprite[0][55][49] = 1;dino_sprite[0][55][50] = 1;dino_sprite[0][55][51] = 1;dino_sprite[0][55][52] = 1;dino_sprite[0][55][53] = 1;dino_sprite[0][55][54] = 1;dino_sprite[0][55][55] = 1;dino_sprite[0][55][56] = 1;dino_sprite[0][55][57] = 1;dino_sprite[0][55][58] = 1;dino_sprite[0][55][59] = 1;dino_sprite[0][55][60] = 1;dino_sprite[0][55][61] = 1;dino_sprite[0][55][62] = 1;dino_sprite[0][55][63] = 1;dino_sprite[0][55][64] = 1;dino_sprite[0][55][65] = 1;dino_sprite[0][55][66] = 1;dino_sprite[0][55][67] = 1;dino_sprite[0][55][68] = 1;dino_sprite[0][55][69] = 1;dino_sprite[0][55][70] = 1;dino_sprite[0][55][71] = 1;dino_sprite[0][55][72] = 1;dino_sprite[0][55][73] = 1;dino_sprite[0][55][74] = 1;dino_sprite[0][55][75] = 1;dino_sprite[0][55][76] = 1;dino_sprite[0][55][77] = 1;dino_sprite[0][55][78] = 1;dino_sprite[0][55][79] = 1;dino_sprite[0][55][80] = 1;dino_sprite[0][55][81] = 1;dino_sprite[0][55][82] = 1;dino_sprite[0][55][83] = 1;dino_sprite[0][55][84] = 1;dino_sprite[0][55][85] = 1;dino_sprite[0][55][86] = 1;dino_sprite[0][55][87] = 1;dino_sprite[0][55][88] = 1;dino_sprite[0][55][89] = 1;dino_sprite[0][55][90] = 1;dino_sprite[0][55][91] = 1;dino_sprite[0][55][92] = 1;dino_sprite[0][55][93] = 1;dino_sprite[0][55][94] = 1;dino_sprite[0][55][95] = 1;dino_sprite[0][55][96] = 1;dino_sprite[0][55][97] = 1;dino_sprite[0][55][98] = 1;dino_sprite[0][55][99] = 1;dino_sprite[0][56][0] = 1;dino_sprite[0][56][1] = 1;dino_sprite[0][56][2] = 1;dino_sprite[0][56][3] = 1;dino_sprite[0][56][4] = 1;dino_sprite[0][56][5] = 1;dino_sprite[0][56][6] = 1;dino_sprite[0][56][7] = 1;dino_sprite[0][56][8] = 1;dino_sprite[0][56][9] = 1;dino_sprite[0][56][10] = 1;dino_sprite[0][56][11] = 1;dino_sprite[0][56][12] = 1;dino_sprite[0][56][13] = 1;dino_sprite[0][56][14] = 1;dino_sprite[0][56][15] = 1;dino_sprite[0][56][16] = 1;dino_sprite[0][56][17] = 1;dino_sprite[0][56][18] = 1;dino_sprite[0][56][19] = 1;dino_sprite[0][56][20] = 1;dino_sprite[0][56][21] = 1;dino_sprite[0][56][22] = 1;dino_sprite[0][56][23] = 1;dino_sprite[0][56][24] = 1;dino_sprite[0][56][25] = 1;dino_sprite[0][56][26] = 1;dino_sprite[0][56][27] = 1;dino_sprite[0][56][28] = 1;dino_sprite[0][56][29] = 1;dino_sprite[0][56][30] = 1;dino_sprite[0][56][31] = 1;dino_sprite[0][56][32] = 1;dino_sprite[0][56][33] = 1;dino_sprite[0][56][34] = 1;dino_sprite[0][56][35] = 1;dino_sprite[0][56][36] = 1;dino_sprite[0][56][37] = 1;dino_sprite[0][56][38] = 1;dino_sprite[0][56][39] = 1;dino_sprite[0][56][40] = 1;dino_sprite[0][56][41] = 1;dino_sprite[0][56][42] = 1;dino_sprite[0][56][43] = 1;dino_sprite[0][56][44] = 1;dino_sprite[0][56][45] = 1;dino_sprite[0][56][46] = 1;dino_sprite[0][56][47] = 1;dino_sprite[0][56][48] = 1;dino_sprite[0][56][49] = 1;dino_sprite[0][56][50] = 1;dino_sprite[0][56][51] = 1;dino_sprite[0][56][52] = 1;dino_sprite[0][56][53] = 1;dino_sprite[0][56][54] = 1;dino_sprite[0][56][55] = 1;dino_sprite[0][56][56] = 1;dino_sprite[0][56][57] = 1;dino_sprite[0][56][58] = 1;dino_sprite[0][56][59] = 1;dino_sprite[0][56][60] = 1;dino_sprite[0][56][61] = 1;dino_sprite[0][56][62] = 1;dino_sprite[0][56][63] = 1;dino_sprite[0][56][64] = 1;dino_sprite[0][56][65] = 1;dino_sprite[0][56][66] = 1;dino_sprite[0][56][67] = 1;dino_sprite[0][56][68] = 1;dino_sprite[0][56][69] = 1;dino_sprite[0][56][70] = 1;dino_sprite[0][56][71] = 1;dino_sprite[0][56][72] = 1;dino_sprite[0][56][73] = 1;dino_sprite[0][56][74] = 1;dino_sprite[0][56][75] = 1;dino_sprite[0][56][76] = 1;dino_sprite[0][56][77] = 1;dino_sprite[0][56][95] = 1;dino_sprite[0][56][96] = 1;dino_sprite[0][56][97] = 1;dino_sprite[0][56][98] = 1;dino_sprite[0][56][99] = 1;dino_sprite[0][57][0] = 1;dino_sprite[0][57][1] = 1;dino_sprite[0][57][2] = 1;dino_sprite[0][57][3] = 1;dino_sprite[0][57][4] = 1;dino_sprite[0][57][5] = 1;dino_sprite[0][57][6] = 1;dino_sprite[0][57][7] = 1;dino_sprite[0][57][8] = 1;dino_sprite[0][57][9] = 1;dino_sprite[0][57][10] = 1;dino_sprite[0][57][11] = 1;dino_sprite[0][57][12] = 1;dino_sprite[0][57][13] = 1;dino_sprite[0][57][14] = 1;dino_sprite[0][57][15] = 1;dino_sprite[0][57][16] = 1;dino_sprite[0][57][17] = 1;dino_sprite[0][57][18] = 1;dino_sprite[0][57][19] = 1;dino_sprite[0][57][20] = 1;dino_sprite[0][57][21] = 1;dino_sprite[0][57][22] = 1;dino_sprite[0][57][23] = 1;dino_sprite[0][57][24] = 1;dino_sprite[0][57][25] = 1;dino_sprite[0][57][26] = 1;dino_sprite[0][57][27] = 1;dino_sprite[0][57][28] = 1;dino_sprite[0][57][29] = 1;dino_sprite[0][57][30] = 1;dino_sprite[0][57][31] = 1;dino_sprite[0][57][32] = 1;dino_sprite[0][57][33] = 1;dino_sprite[0][57][34] = 1;dino_sprite[0][57][35] = 1;dino_sprite[0][57][36] = 1;dino_sprite[0][57][37] = 1;dino_sprite[0][57][38] = 1;dino_sprite[0][57][39] = 1;dino_sprite[0][57][40] = 1;dino_sprite[0][57][41] = 1;dino_sprite[0][57][42] = 1;dino_sprite[0][57][43] = 1;dino_sprite[0][57][44] = 1;dino_sprite[0][57][45] = 1;dino_sprite[0][57][46] = 1;dino_sprite[0][57][47] = 1;dino_sprite[0][57][48] = 1;dino_sprite[0][57][49] = 1;dino_sprite[0][57][50] = 1;dino_sprite[0][57][51] = 1;dino_sprite[0][57][52] = 1;dino_sprite[0][57][53] = 1;dino_sprite[0][57][54] = 1;dino_sprite[0][57][55] = 1;dino_sprite[0][57][56] = 1;dino_sprite[0][57][57] = 1;dino_sprite[0][57][58] = 1;dino_sprite[0][57][59] = 1;dino_sprite[0][57][60] = 1;dino_sprite[0][57][61] = 1;dino_sprite[0][57][62] = 1;dino_sprite[0][57][63] = 1;dino_sprite[0][57][64] = 1;dino_sprite[0][57][65] = 1;dino_sprite[0][57][66] = 1;dino_sprite[0][57][67] = 1;dino_sprite[0][57][68] = 1;dino_sprite[0][57][69] = 1;dino_sprite[0][57][70] = 1;dino_sprite[0][57][71] = 1;dino_sprite[0][57][72] = 1;dino_sprite[0][57][73] = 1;dino_sprite[0][57][74] = 1;dino_sprite[0][57][75] = 1;dino_sprite[0][57][76] = 1;dino_sprite[0][57][77] = 1;dino_sprite[0][57][95] = 1;dino_sprite[0][57][96] = 1;dino_sprite[0][57][97] = 1;dino_sprite[0][57][98] = 1;dino_sprite[0][57][99] = 1;dino_sprite[0][58][0] = 1;dino_sprite[0][58][1] = 1;dino_sprite[0][58][2] = 1;dino_sprite[0][58][3] = 1;dino_sprite[0][58][4] = 1;dino_sprite[0][58][5] = 1;dino_sprite[0][58][6] = 1;dino_sprite[0][58][7] = 1;dino_sprite[0][58][8] = 1;dino_sprite[0][58][9] = 1;dino_sprite[0][58][10] = 1;dino_sprite[0][58][11] = 1;dino_sprite[0][58][12] = 1;dino_sprite[0][58][13] = 1;dino_sprite[0][58][14] = 1;dino_sprite[0][58][15] = 1;dino_sprite[0][58][16] = 1;dino_sprite[0][58][17] = 1;dino_sprite[0][58][18] = 1;dino_sprite[0][58][19] = 1;dino_sprite[0][58][20] = 1;dino_sprite[0][58][21] = 1;dino_sprite[0][58][22] = 1;dino_sprite[0][58][23] = 1;dino_sprite[0][58][24] = 1;dino_sprite[0][58][25] = 1;dino_sprite[0][58][26] = 1;dino_sprite[0][58][27] = 1;dino_sprite[0][58][28] = 1;dino_sprite[0][58][29] = 1;dino_sprite[0][58][30] = 1;dino_sprite[0][58][31] = 1;dino_sprite[0][58][32] = 1;dino_sprite[0][58][33] = 1;dino_sprite[0][58][34] = 1;dino_sprite[0][58][35] = 1;dino_sprite[0][58][36] = 1;dino_sprite[0][58][37] = 1;dino_sprite[0][58][38] = 1;dino_sprite[0][58][39] = 1;dino_sprite[0][58][40] = 1;dino_sprite[0][58][41] = 1;dino_sprite[0][58][42] = 1;dino_sprite[0][58][43] = 1;dino_sprite[0][58][44] = 1;dino_sprite[0][58][45] = 1;dino_sprite[0][58][46] = 1;dino_sprite[0][58][47] = 1;dino_sprite[0][58][48] = 1;dino_sprite[0][58][49] = 1;dino_sprite[0][58][50] = 1;dino_sprite[0][58][51] = 1;dino_sprite[0][58][52] = 1;dino_sprite[0][58][53] = 1;dino_sprite[0][58][54] = 1;dino_sprite[0][58][55] = 1;dino_sprite[0][58][56] = 1;dino_sprite[0][58][57] = 1;dino_sprite[0][58][58] = 1;dino_sprite[0][58][59] = 1;dino_sprite[0][58][60] = 1;dino_sprite[0][58][61] = 1;dino_sprite[0][58][62] = 1;dino_sprite[0][58][63] = 1;dino_sprite[0][58][64] = 1;dino_sprite[0][58][65] = 1;dino_sprite[0][58][66] = 1;dino_sprite[0][58][67] = 1;dino_sprite[0][58][68] = 1;dino_sprite[0][58][69] = 1;dino_sprite[0][58][70] = 1;dino_sprite[0][58][71] = 1;dino_sprite[0][58][72] = 1;dino_sprite[0][58][73] = 1;dino_sprite[0][58][74] = 1;dino_sprite[0][58][75] = 1;dino_sprite[0][58][76] = 1;dino_sprite[0][58][77] = 1;dino_sprite[0][58][95] = 1;dino_sprite[0][58][96] = 1;dino_sprite[0][58][97] = 1;dino_sprite[0][58][98] = 1;dino_sprite[0][58][99] = 1;dino_sprite[0][59][0] = 1;dino_sprite[0][59][1] = 1;dino_sprite[0][59][2] = 1;dino_sprite[0][59][3] = 1;dino_sprite[0][59][4] = 1;dino_sprite[0][59][5] = 1;dino_sprite[0][59][6] = 1;dino_sprite[0][59][7] = 1;dino_sprite[0][59][8] = 1;dino_sprite[0][59][9] = 1;dino_sprite[0][59][10] = 1;dino_sprite[0][59][11] = 1;dino_sprite[0][59][12] = 1;dino_sprite[0][59][13] = 1;dino_sprite[0][59][14] = 1;dino_sprite[0][59][15] = 1;dino_sprite[0][59][16] = 1;dino_sprite[0][59][17] = 1;dino_sprite[0][59][18] = 1;dino_sprite[0][59][19] = 1;dino_sprite[0][59][20] = 1;dino_sprite[0][59][21] = 1;dino_sprite[0][59][22] = 1;dino_sprite[0][59][23] = 1;dino_sprite[0][59][24] = 1;dino_sprite[0][59][25] = 1;dino_sprite[0][59][26] = 1;dino_sprite[0][59][27] = 1;dino_sprite[0][59][28] = 1;dino_sprite[0][59][29] = 1;dino_sprite[0][59][30] = 1;dino_sprite[0][59][31] = 1;dino_sprite[0][59][32] = 1;dino_sprite[0][59][33] = 1;dino_sprite[0][59][34] = 1;dino_sprite[0][59][35] = 1;dino_sprite[0][59][36] = 1;dino_sprite[0][59][37] = 1;dino_sprite[0][59][38] = 1;dino_sprite[0][59][39] = 1;dino_sprite[0][59][40] = 1;dino_sprite[0][59][41] = 1;dino_sprite[0][59][42] = 1;dino_sprite[0][59][43] = 1;dino_sprite[0][59][44] = 1;dino_sprite[0][59][45] = 1;dino_sprite[0][59][46] = 1;dino_sprite[0][59][47] = 1;dino_sprite[0][59][48] = 1;dino_sprite[0][59][49] = 1;dino_sprite[0][59][50] = 1;dino_sprite[0][59][51] = 1;dino_sprite[0][59][52] = 1;dino_sprite[0][59][53] = 1;dino_sprite[0][59][54] = 1;dino_sprite[0][59][55] = 1;dino_sprite[0][59][56] = 1;dino_sprite[0][59][57] = 1;dino_sprite[0][59][58] = 1;dino_sprite[0][59][59] = 1;dino_sprite[0][59][60] = 1;dino_sprite[0][59][61] = 1;dino_sprite[0][59][62] = 1;dino_sprite[0][59][63] = 1;dino_sprite[0][59][64] = 1;dino_sprite[0][59][65] = 1;dino_sprite[0][59][66] = 1;dino_sprite[0][59][67] = 1;dino_sprite[0][59][68] = 1;dino_sprite[0][59][69] = 1;dino_sprite[0][59][70] = 1;dino_sprite[0][59][71] = 1;dino_sprite[0][59][72] = 1;dino_sprite[0][59][73] = 1;dino_sprite[0][59][74] = 1;dino_sprite[0][59][75] = 1;dino_sprite[0][59][76] = 1;dino_sprite[0][59][77] = 1;dino_sprite[0][59][95] = 1;dino_sprite[0][59][96] = 1;dino_sprite[0][59][97] = 1;dino_sprite[0][59][98] = 1;dino_sprite[0][59][99] = 1;dino_sprite[0][60][0] = 1;dino_sprite[0][60][1] = 1;dino_sprite[0][60][2] = 1;dino_sprite[0][60][3] = 1;dino_sprite[0][60][4] = 1;dino_sprite[0][60][5] = 1;dino_sprite[0][60][6] = 1;dino_sprite[0][60][7] = 1;dino_sprite[0][60][8] = 1;dino_sprite[0][60][9] = 1;dino_sprite[0][60][10] = 1;dino_sprite[0][60][11] = 1;dino_sprite[0][60][12] = 1;dino_sprite[0][60][13] = 1;dino_sprite[0][60][14] = 1;dino_sprite[0][60][15] = 1;dino_sprite[0][60][16] = 1;dino_sprite[0][60][17] = 1;dino_sprite[0][60][18] = 1;dino_sprite[0][60][19] = 1;dino_sprite[0][60][20] = 1;dino_sprite[0][60][21] = 1;dino_sprite[0][60][22] = 1;dino_sprite[0][60][23] = 1;dino_sprite[0][60][24] = 1;dino_sprite[0][60][25] = 1;dino_sprite[0][60][26] = 1;dino_sprite[0][60][27] = 1;dino_sprite[0][60][28] = 1;dino_sprite[0][60][29] = 1;dino_sprite[0][60][30] = 1;dino_sprite[0][60][31] = 1;dino_sprite[0][60][32] = 1;dino_sprite[0][60][33] = 1;dino_sprite[0][60][34] = 1;dino_sprite[0][60][35] = 1;dino_sprite[0][60][36] = 1;dino_sprite[0][60][37] = 1;dino_sprite[0][60][38] = 1;dino_sprite[0][60][39] = 1;dino_sprite[0][60][40] = 1;dino_sprite[0][60][41] = 1;dino_sprite[0][60][42] = 1;dino_sprite[0][60][43] = 1;dino_sprite[0][60][44] = 1;dino_sprite[0][60][45] = 1;dino_sprite[0][60][46] = 1;dino_sprite[0][60][47] = 1;dino_sprite[0][60][48] = 1;dino_sprite[0][60][49] = 1;dino_sprite[0][60][50] = 1;dino_sprite[0][60][51] = 1;dino_sprite[0][60][52] = 1;dino_sprite[0][60][53] = 1;dino_sprite[0][60][54] = 1;dino_sprite[0][60][55] = 1;dino_sprite[0][60][56] = 1;dino_sprite[0][60][57] = 1;dino_sprite[0][60][58] = 1;dino_sprite[0][60][59] = 1;dino_sprite[0][60][60] = 1;dino_sprite[0][60][61] = 1;dino_sprite[0][60][62] = 1;dino_sprite[0][60][63] = 1;dino_sprite[0][60][64] = 1;dino_sprite[0][60][65] = 1;dino_sprite[0][60][66] = 1;dino_sprite[0][60][67] = 1;dino_sprite[0][60][68] = 1;dino_sprite[0][60][69] = 1;dino_sprite[0][60][70] = 1;dino_sprite[0][60][71] = 1;dino_sprite[0][60][72] = 1;dino_sprite[0][60][73] = 1;dino_sprite[0][60][74] = 1;dino_sprite[0][60][75] = 1;dino_sprite[0][60][76] = 1;dino_sprite[0][60][77] = 1;dino_sprite[0][60][96] = 1;dino_sprite[0][60][97] = 1;dino_sprite[0][60][98] = 1;dino_sprite[0][60][99] = 1;dino_sprite[0][61][0] = 1;dino_sprite[0][61][1] = 1;dino_sprite[0][61][2] = 1;dino_sprite[0][61][3] = 1;dino_sprite[0][61][4] = 1;dino_sprite[0][61][5] = 1;dino_sprite[0][61][6] = 1;dino_sprite[0][61][10] = 1;dino_sprite[0][61][11] = 1;dino_sprite[0][61][12] = 1;dino_sprite[0][61][13] = 1;dino_sprite[0][61][14] = 1;dino_sprite[0][61][15] = 1;dino_sprite[0][61][16] = 1;dino_sprite[0][61][17] = 1;dino_sprite[0][61][18] = 1;dino_sprite[0][61][19] = 1;dino_sprite[0][61][20] = 1;dino_sprite[0][61][21] = 1;dino_sprite[0][61][22] = 1;dino_sprite[0][61][23] = 1;dino_sprite[0][61][24] = 1;dino_sprite[0][61][25] = 1;dino_sprite[0][61][26] = 1;dino_sprite[0][61][27] = 1;dino_sprite[0][61][28] = 1;dino_sprite[0][61][29] = 1;dino_sprite[0][61][30] = 1;dino_sprite[0][61][31] = 1;dino_sprite[0][61][32] = 1;dino_sprite[0][61][33] = 1;dino_sprite[0][61][34] = 1;dino_sprite[0][61][35] = 1;dino_sprite[0][61][36] = 1;dino_sprite[0][61][37] = 1;dino_sprite[0][61][38] = 1;dino_sprite[0][61][39] = 1;dino_sprite[0][61][40] = 1;dino_sprite[0][61][41] = 1;dino_sprite[0][61][42] = 1;dino_sprite[0][61][43] = 1;dino_sprite[0][61][44] = 1;dino_sprite[0][61][45] = 1;dino_sprite[0][61][46] = 1;dino_sprite[0][61][47] = 1;dino_sprite[0][61][48] = 1;dino_sprite[0][61][49] = 1;dino_sprite[0][61][50] = 1;dino_sprite[0][61][51] = 1;dino_sprite[0][61][52] = 1;dino_sprite[0][61][53] = 1;dino_sprite[0][61][54] = 1;dino_sprite[0][61][55] = 1;dino_sprite[0][61][56] = 1;dino_sprite[0][61][57] = 1;dino_sprite[0][61][58] = 1;dino_sprite[0][61][59] = 1;dino_sprite[0][61][60] = 1;dino_sprite[0][61][61] = 1;dino_sprite[0][61][62] = 1;dino_sprite[0][61][63] = 1;dino_sprite[0][61][64] = 1;dino_sprite[0][61][65] = 1;dino_sprite[0][61][66] = 1;dino_sprite[0][61][67] = 1;dino_sprite[0][61][68] = 1;dino_sprite[0][61][69] = 1;dino_sprite[0][61][70] = 1;dino_sprite[0][61][71] = 1;dino_sprite[0][61][72] = 1;dino_sprite[0][62][0] = 1;dino_sprite[0][62][1] = 1;dino_sprite[0][62][2] = 1;dino_sprite[0][62][3] = 1;dino_sprite[0][62][4] = 1;dino_sprite[0][62][5] = 1;dino_sprite[0][62][6] = 1;dino_sprite[0][62][10] = 1;dino_sprite[0][62][11] = 1;dino_sprite[0][62][12] = 1;dino_sprite[0][62][13] = 1;dino_sprite[0][62][14] = 1;dino_sprite[0][62][15] = 1;dino_sprite[0][62][16] = 1;dino_sprite[0][62][17] = 1;dino_sprite[0][62][18] = 1;dino_sprite[0][62][19] = 1;dino_sprite[0][62][20] = 1;dino_sprite[0][62][21] = 1;dino_sprite[0][62][22] = 1;dino_sprite[0][62][23] = 1;dino_sprite[0][62][24] = 1;dino_sprite[0][62][25] = 1;dino_sprite[0][62][26] = 1;dino_sprite[0][62][27] = 1;dino_sprite[0][62][28] = 1;dino_sprite[0][62][29] = 1;dino_sprite[0][62][30] = 1;dino_sprite[0][62][31] = 1;dino_sprite[0][62][32] = 1;dino_sprite[0][62][33] = 1;dino_sprite[0][62][34] = 1;dino_sprite[0][62][35] = 1;dino_sprite[0][62][36] = 1;dino_sprite[0][62][37] = 1;dino_sprite[0][62][38] = 1;dino_sprite[0][62][39] = 1;dino_sprite[0][62][40] = 1;dino_sprite[0][62][41] = 1;dino_sprite[0][62][42] = 1;dino_sprite[0][62][43] = 1;dino_sprite[0][62][44] = 1;dino_sprite[0][62][45] = 1;dino_sprite[0][62][46] = 1;dino_sprite[0][62][47] = 1;dino_sprite[0][62][48] = 1;dino_sprite[0][62][49] = 1;dino_sprite[0][62][50] = 1;dino_sprite[0][62][51] = 1;dino_sprite[0][62][52] = 1;dino_sprite[0][62][53] = 1;dino_sprite[0][62][54] = 1;dino_sprite[0][62][55] = 1;dino_sprite[0][62][56] = 1;dino_sprite[0][62][57] = 1;dino_sprite[0][62][58] = 1;dino_sprite[0][62][59] = 1;dino_sprite[0][62][60] = 1;dino_sprite[0][62][61] = 1;dino_sprite[0][62][62] = 1;dino_sprite[0][62][63] = 1;dino_sprite[0][62][64] = 1;dino_sprite[0][62][65] = 1;dino_sprite[0][62][66] = 1;dino_sprite[0][62][67] = 1;dino_sprite[0][62][68] = 1;dino_sprite[0][62][69] = 1;dino_sprite[0][62][70] = 1;dino_sprite[0][62][71] = 1;dino_sprite[0][62][72] = 1;dino_sprite[0][63][0] = 1;dino_sprite[0][63][1] = 1;dino_sprite[0][63][2] = 1;dino_sprite[0][63][3] = 1;dino_sprite[0][63][4] = 1;dino_sprite[0][63][5] = 1;dino_sprite[0][63][6] = 1;dino_sprite[0][63][10] = 1;dino_sprite[0][63][11] = 1;dino_sprite[0][63][12] = 1;dino_sprite[0][63][13] = 1;dino_sprite[0][63][14] = 1;dino_sprite[0][63][15] = 1;dino_sprite[0][63][16] = 1;dino_sprite[0][63][17] = 1;dino_sprite[0][63][18] = 1;dino_sprite[0][63][19] = 1;dino_sprite[0][63][20] = 1;dino_sprite[0][63][21] = 1;dino_sprite[0][63][22] = 1;dino_sprite[0][63][23] = 1;dino_sprite[0][63][24] = 1;dino_sprite[0][63][25] = 1;dino_sprite[0][63][26] = 1;dino_sprite[0][63][27] = 1;dino_sprite[0][63][28] = 1;dino_sprite[0][63][29] = 1;dino_sprite[0][63][30] = 1;dino_sprite[0][63][31] = 1;dino_sprite[0][63][32] = 1;dino_sprite[0][63][33] = 1;dino_sprite[0][63][34] = 1;dino_sprite[0][63][35] = 1;dino_sprite[0][63][36] = 1;dino_sprite[0][63][37] = 1;dino_sprite[0][63][38] = 1;dino_sprite[0][63][39] = 1;dino_sprite[0][63][40] = 1;dino_sprite[0][63][41] = 1;dino_sprite[0][63][42] = 1;dino_sprite[0][63][43] = 1;dino_sprite[0][63][44] = 1;dino_sprite[0][63][45] = 1;dino_sprite[0][63][46] = 1;dino_sprite[0][63][47] = 1;dino_sprite[0][63][48] = 1;dino_sprite[0][63][49] = 1;dino_sprite[0][63][50] = 1;dino_sprite[0][63][51] = 1;dino_sprite[0][63][52] = 1;dino_sprite[0][63][53] = 1;dino_sprite[0][63][54] = 1;dino_sprite[0][63][55] = 1;dino_sprite[0][63][56] = 1;dino_sprite[0][63][57] = 1;dino_sprite[0][63][58] = 1;dino_sprite[0][63][59] = 1;dino_sprite[0][63][60] = 1;dino_sprite[0][63][61] = 1;dino_sprite[0][63][62] = 1;dino_sprite[0][63][63] = 1;dino_sprite[0][63][64] = 1;dino_sprite[0][63][65] = 1;dino_sprite[0][63][66] = 1;dino_sprite[0][63][67] = 1;dino_sprite[0][63][68] = 1;dino_sprite[0][63][69] = 1;dino_sprite[0][63][70] = 1;dino_sprite[0][63][71] = 1;dino_sprite[0][63][72] = 1;dino_sprite[0][64][0] = 1;dino_sprite[0][64][1] = 1;dino_sprite[0][64][2] = 1;dino_sprite[0][64][3] = 1;dino_sprite[0][64][4] = 1;dino_sprite[0][64][5] = 1;dino_sprite[0][64][6] = 1;dino_sprite[0][64][10] = 1;dino_sprite[0][64][11] = 1;dino_sprite[0][64][12] = 1;dino_sprite[0][64][13] = 1;dino_sprite[0][64][14] = 1;dino_sprite[0][64][15] = 1;dino_sprite[0][64][16] = 1;dino_sprite[0][64][17] = 1;dino_sprite[0][64][18] = 1;dino_sprite[0][64][19] = 1;dino_sprite[0][64][20] = 1;dino_sprite[0][64][21] = 1;dino_sprite[0][64][22] = 1;dino_sprite[0][64][23] = 1;dino_sprite[0][64][24] = 1;dino_sprite[0][64][25] = 1;dino_sprite[0][64][26] = 1;dino_sprite[0][64][27] = 1;dino_sprite[0][64][28] = 1;dino_sprite[0][64][29] = 1;dino_sprite[0][64][30] = 1;dino_sprite[0][64][31] = 1;dino_sprite[0][64][32] = 1;dino_sprite[0][64][33] = 1;dino_sprite[0][64][34] = 1;dino_sprite[0][64][35] = 1;dino_sprite[0][64][36] = 1;dino_sprite[0][64][37] = 1;dino_sprite[0][64][38] = 1;dino_sprite[0][64][39] = 1;dino_sprite[0][64][40] = 1;dino_sprite[0][64][41] = 1;dino_sprite[0][64][42] = 1;dino_sprite[0][64][43] = 1;dino_sprite[0][64][44] = 1;dino_sprite[0][64][45] = 1;dino_sprite[0][64][46] = 1;dino_sprite[0][64][47] = 1;dino_sprite[0][64][48] = 1;dino_sprite[0][64][49] = 1;dino_sprite[0][64][50] = 1;dino_sprite[0][64][51] = 1;dino_sprite[0][64][52] = 1;dino_sprite[0][64][53] = 1;dino_sprite[0][64][54] = 1;dino_sprite[0][64][55] = 1;dino_sprite[0][64][56] = 1;dino_sprite[0][64][57] = 1;dino_sprite[0][64][58] = 1;dino_sprite[0][64][59] = 1;dino_sprite[0][64][60] = 1;dino_sprite[0][64][61] = 1;dino_sprite[0][64][62] = 1;dino_sprite[0][64][63] = 1;dino_sprite[0][64][64] = 1;dino_sprite[0][64][65] = 1;dino_sprite[0][64][66] = 1;dino_sprite[0][64][67] = 1;dino_sprite[0][64][68] = 1;dino_sprite[0][64][69] = 1;dino_sprite[0][64][70] = 1;dino_sprite[0][64][71] = 1;dino_sprite[0][64][72] = 1;dino_sprite[0][65][0] = 1;dino_sprite[0][65][1] = 1;dino_sprite[0][65][2] = 1;dino_sprite[0][65][3] = 1;dino_sprite[0][65][4] = 1;dino_sprite[0][65][5] = 1;dino_sprite[0][65][6] = 1;dino_sprite[0][65][8] = 1;dino_sprite[0][65][10] = 1;dino_sprite[0][65][11] = 1;dino_sprite[0][65][12] = 1;dino_sprite[0][65][13] = 1;dino_sprite[0][65][14] = 1;dino_sprite[0][65][15] = 1;dino_sprite[0][65][16] = 1;dino_sprite[0][65][17] = 1;dino_sprite[0][65][18] = 1;dino_sprite[0][65][19] = 1;dino_sprite[0][65][20] = 1;dino_sprite[0][65][21] = 1;dino_sprite[0][65][22] = 1;dino_sprite[0][65][23] = 1;dino_sprite[0][65][24] = 1;dino_sprite[0][65][25] = 1;dino_sprite[0][65][26] = 1;dino_sprite[0][65][27] = 1;dino_sprite[0][65][28] = 1;dino_sprite[0][65][29] = 1;dino_sprite[0][65][30] = 1;dino_sprite[0][65][31] = 1;dino_sprite[0][65][32] = 1;dino_sprite[0][65][33] = 1;dino_sprite[0][65][34] = 1;dino_sprite[0][65][35] = 1;dino_sprite[0][65][36] = 1;dino_sprite[0][65][37] = 1;dino_sprite[0][65][38] = 1;dino_sprite[0][65][39] = 1;dino_sprite[0][65][40] = 1;dino_sprite[0][65][41] = 1;dino_sprite[0][65][42] = 1;dino_sprite[0][65][43] = 1;dino_sprite[0][65][44] = 1;dino_sprite[0][65][45] = 1;dino_sprite[0][65][46] = 1;dino_sprite[0][65][47] = 1;dino_sprite[0][65][48] = 1;dino_sprite[0][65][49] = 1;dino_sprite[0][65][50] = 1;dino_sprite[0][65][51] = 1;dino_sprite[0][65][52] = 1;dino_sprite[0][65][53] = 1;dino_sprite[0][65][54] = 1;dino_sprite[0][65][55] = 1;dino_sprite[0][65][56] = 1;dino_sprite[0][65][57] = 1;dino_sprite[0][65][58] = 1;dino_sprite[0][65][59] = 1;dino_sprite[0][65][60] = 1;dino_sprite[0][65][61] = 1;dino_sprite[0][65][62] = 1;dino_sprite[0][65][63] = 1;dino_sprite[0][65][64] = 1;dino_sprite[0][65][65] = 1;dino_sprite[0][65][66] = 1;dino_sprite[0][65][67] = 1;dino_sprite[0][65][68] = 1;dino_sprite[0][65][69] = 1;dino_sprite[0][65][70] = 1;dino_sprite[0][65][71] = 1;dino_sprite[0][65][72] = 1;dino_sprite[0][66][0] = 1;dino_sprite[0][66][1] = 1;dino_sprite[0][66][2] = 1;dino_sprite[0][66][3] = 1;dino_sprite[0][66][4] = 1;dino_sprite[0][66][5] = 1;dino_sprite[0][66][6] = 1;dino_sprite[0][66][7] = 1;dino_sprite[0][66][8] = 1;dino_sprite[0][66][9] = 1;dino_sprite[0][66][10] = 1;dino_sprite[0][66][11] = 1;dino_sprite[0][66][12] = 1;dino_sprite[0][66][13] = 1;dino_sprite[0][66][14] = 1;dino_sprite[0][66][15] = 1;dino_sprite[0][66][16] = 1;dino_sprite[0][66][17] = 1;dino_sprite[0][66][18] = 1;dino_sprite[0][66][19] = 1;dino_sprite[0][66][20] = 1;dino_sprite[0][66][21] = 1;dino_sprite[0][66][22] = 1;dino_sprite[0][66][23] = 1;dino_sprite[0][66][24] = 1;dino_sprite[0][66][25] = 1;dino_sprite[0][66][26] = 1;dino_sprite[0][66][27] = 1;dino_sprite[0][66][28] = 1;dino_sprite[0][66][29] = 1;dino_sprite[0][66][30] = 1;dino_sprite[0][66][31] = 1;dino_sprite[0][66][32] = 1;dino_sprite[0][66][33] = 1;dino_sprite[0][66][34] = 1;dino_sprite[0][66][35] = 1;dino_sprite[0][66][36] = 1;dino_sprite[0][66][37] = 1;dino_sprite[0][66][38] = 1;dino_sprite[0][66][39] = 1;dino_sprite[0][66][40] = 1;dino_sprite[0][66][41] = 1;dino_sprite[0][66][42] = 1;dino_sprite[0][66][43] = 1;dino_sprite[0][66][44] = 1;dino_sprite[0][66][45] = 1;dino_sprite[0][66][46] = 1;dino_sprite[0][66][47] = 1;dino_sprite[0][66][48] = 1;dino_sprite[0][66][49] = 1;dino_sprite[0][66][50] = 1;dino_sprite[0][66][51] = 1;dino_sprite[0][66][52] = 1;dino_sprite[0][66][53] = 1;dino_sprite[0][66][54] = 1;dino_sprite[0][66][55] = 1;dino_sprite[0][66][56] = 1;dino_sprite[0][66][57] = 1;dino_sprite[0][66][58] = 1;dino_sprite[0][66][59] = 1;dino_sprite[0][66][60] = 1;dino_sprite[0][66][61] = 1;dino_sprite[0][66][62] = 1;dino_sprite[0][66][63] = 1;dino_sprite[0][66][64] = 1;dino_sprite[0][66][65] = 1;dino_sprite[0][67][0] = 1;dino_sprite[0][67][1] = 1;dino_sprite[0][67][2] = 1;dino_sprite[0][67][3] = 1;dino_sprite[0][67][4] = 1;dino_sprite[0][67][5] = 1;dino_sprite[0][67][6] = 1;dino_sprite[0][67][7] = 1;dino_sprite[0][67][8] = 1;dino_sprite[0][67][9] = 1;dino_sprite[0][67][10] = 1;dino_sprite[0][67][11] = 1;dino_sprite[0][67][12] = 1;dino_sprite[0][67][13] = 1;dino_sprite[0][67][14] = 1;dino_sprite[0][67][15] = 1;dino_sprite[0][67][16] = 1;dino_sprite[0][67][17] = 1;dino_sprite[0][67][18] = 1;dino_sprite[0][67][19] = 1;dino_sprite[0][67][20] = 1;dino_sprite[0][67][21] = 1;dino_sprite[0][67][22] = 1;dino_sprite[0][67][23] = 1;dino_sprite[0][67][24] = 1;dino_sprite[0][67][25] = 1;dino_sprite[0][67][26] = 1;dino_sprite[0][67][27] = 1;dino_sprite[0][67][28] = 1;dino_sprite[0][67][29] = 1;dino_sprite[0][67][30] = 1;dino_sprite[0][67][31] = 1;dino_sprite[0][67][32] = 1;dino_sprite[0][67][33] = 1;dino_sprite[0][67][34] = 1;dino_sprite[0][67][35] = 1;dino_sprite[0][67][36] = 1;dino_sprite[0][67][37] = 1;dino_sprite[0][67][38] = 1;dino_sprite[0][67][39] = 1;dino_sprite[0][67][40] = 1;dino_sprite[0][67][41] = 1;dino_sprite[0][67][42] = 1;dino_sprite[0][67][43] = 1;dino_sprite[0][67][44] = 1;dino_sprite[0][67][45] = 1;dino_sprite[0][67][46] = 1;dino_sprite[0][67][47] = 1;dino_sprite[0][67][48] = 1;dino_sprite[0][67][49] = 1;dino_sprite[0][67][50] = 1;dino_sprite[0][67][51] = 1;dino_sprite[0][67][52] = 1;dino_sprite[0][67][53] = 1;dino_sprite[0][67][54] = 1;dino_sprite[0][67][55] = 1;dino_sprite[0][67][56] = 1;dino_sprite[0][67][57] = 1;dino_sprite[0][67][58] = 1;dino_sprite[0][67][59] = 1;dino_sprite[0][67][60] = 1;dino_sprite[0][67][61] = 1;dino_sprite[0][67][62] = 1;dino_sprite[0][67][63] = 1;dino_sprite[0][67][64] = 1;dino_sprite[0][67][65] = 1;dino_sprite[0][68][0] = 1;dino_sprite[0][68][1] = 1;dino_sprite[0][68][2] = 1;dino_sprite[0][68][3] = 1;dino_sprite[0][68][4] = 1;dino_sprite[0][68][5] = 1;dino_sprite[0][68][6] = 1;dino_sprite[0][68][7] = 1;dino_sprite[0][68][8] = 1;dino_sprite[0][68][9] = 1;dino_sprite[0][68][10] = 1;dino_sprite[0][68][11] = 1;dino_sprite[0][68][12] = 1;dino_sprite[0][68][13] = 1;dino_sprite[0][68][14] = 1;dino_sprite[0][68][15] = 1;dino_sprite[0][68][16] = 1;dino_sprite[0][68][17] = 1;dino_sprite[0][68][18] = 1;dino_sprite[0][68][19] = 1;dino_sprite[0][68][20] = 1;dino_sprite[0][68][21] = 1;dino_sprite[0][68][22] = 1;dino_sprite[0][68][23] = 1;dino_sprite[0][68][24] = 1;dino_sprite[0][68][25] = 1;dino_sprite[0][68][26] = 1;dino_sprite[0][68][27] = 1;dino_sprite[0][68][28] = 1;dino_sprite[0][68][29] = 1;dino_sprite[0][68][30] = 1;dino_sprite[0][68][31] = 1;dino_sprite[0][68][32] = 1;dino_sprite[0][68][33] = 1;dino_sprite[0][68][34] = 1;dino_sprite[0][68][35] = 1;dino_sprite[0][68][36] = 1;dino_sprite[0][68][37] = 1;dino_sprite[0][68][38] = 1;dino_sprite[0][68][39] = 1;dino_sprite[0][68][40] = 1;dino_sprite[0][68][41] = 1;dino_sprite[0][68][42] = 1;dino_sprite[0][68][43] = 1;dino_sprite[0][68][44] = 1;dino_sprite[0][68][45] = 1;dino_sprite[0][68][46] = 1;dino_sprite[0][68][47] = 1;dino_sprite[0][68][48] = 1;dino_sprite[0][68][49] = 1;dino_sprite[0][68][50] = 1;dino_sprite[0][68][51] = 1;dino_sprite[0][68][52] = 1;dino_sprite[0][68][53] = 1;dino_sprite[0][68][54] = 1;dino_sprite[0][68][55] = 1;dino_sprite[0][68][56] = 1;dino_sprite[0][68][57] = 1;dino_sprite[0][68][58] = 1;dino_sprite[0][68][59] = 1;dino_sprite[0][68][60] = 1;dino_sprite[0][68][61] = 1;dino_sprite[0][68][62] = 1;dino_sprite[0][68][63] = 1;dino_sprite[0][68][64] = 1;dino_sprite[0][68][65] = 1;dino_sprite[0][69][0] = 1;dino_sprite[0][69][1] = 1;dino_sprite[0][69][2] = 1;dino_sprite[0][69][3] = 1;dino_sprite[0][69][4] = 1;dino_sprite[0][69][5] = 1;dino_sprite[0][69][6] = 1;dino_sprite[0][69][7] = 1;dino_sprite[0][69][8] = 1;dino_sprite[0][69][9] = 1;dino_sprite[0][69][10] = 1;dino_sprite[0][69][11] = 1;dino_sprite[0][69][12] = 1;dino_sprite[0][69][13] = 1;dino_sprite[0][69][14] = 1;dino_sprite[0][69][15] = 1;dino_sprite[0][69][16] = 1;dino_sprite[0][69][17] = 1;dino_sprite[0][69][18] = 1;dino_sprite[0][69][19] = 1;dino_sprite[0][69][20] = 1;dino_sprite[0][69][21] = 1;dino_sprite[0][69][22] = 1;dino_sprite[0][69][23] = 1;dino_sprite[0][69][24] = 1;dino_sprite[0][69][25] = 1;dino_sprite[0][69][26] = 1;dino_sprite[0][69][27] = 1;dino_sprite[0][69][28] = 1;dino_sprite[0][69][29] = 1;dino_sprite[0][69][30] = 1;dino_sprite[0][69][31] = 1;dino_sprite[0][69][32] = 1;dino_sprite[0][69][33] = 1;dino_sprite[0][69][34] = 1;dino_sprite[0][69][35] = 1;dino_sprite[0][69][36] = 1;dino_sprite[0][69][37] = 1;dino_sprite[0][69][38] = 1;dino_sprite[0][69][39] = 1;dino_sprite[0][69][40] = 1;dino_sprite[0][69][41] = 1;dino_sprite[0][69][42] = 1;dino_sprite[0][69][43] = 1;dino_sprite[0][69][44] = 1;dino_sprite[0][69][45] = 1;dino_sprite[0][69][46] = 1;dino_sprite[0][69][47] = 1;dino_sprite[0][69][48] = 1;dino_sprite[0][69][49] = 1;dino_sprite[0][69][50] = 1;dino_sprite[0][69][51] = 1;dino_sprite[0][69][52] = 1;dino_sprite[0][69][53] = 1;dino_sprite[0][69][54] = 1;dino_sprite[0][69][55] = 1;dino_sprite[0][69][56] = 1;dino_sprite[0][69][57] = 1;dino_sprite[0][69][58] = 1;dino_sprite[0][69][59] = 1;dino_sprite[0][69][60] = 1;dino_sprite[0][69][61] = 1;dino_sprite[0][69][62] = 1;dino_sprite[0][69][63] = 1;dino_sprite[0][69][64] = 1;dino_sprite[0][69][65] = 1;dino_sprite[0][70][0] = 1;dino_sprite[0][70][1] = 1;dino_sprite[0][70][2] = 1;dino_sprite[0][70][3] = 1;dino_sprite[0][70][4] = 1;dino_sprite[0][70][5] = 1;dino_sprite[0][70][6] = 1;dino_sprite[0][70][7] = 1;dino_sprite[0][70][8] = 1;dino_sprite[0][70][9] = 1;dino_sprite[0][70][10] = 1;dino_sprite[0][70][11] = 1;dino_sprite[0][70][12] = 1;dino_sprite[0][70][13] = 1;dino_sprite[0][70][14] = 1;dino_sprite[0][70][15] = 1;dino_sprite[0][70][16] = 1;dino_sprite[0][70][17] = 1;dino_sprite[0][70][18] = 1;dino_sprite[0][70][19] = 1;dino_sprite[0][70][20] = 1;dino_sprite[0][70][21] = 1;dino_sprite[0][70][22] = 1;dino_sprite[0][70][23] = 1;dino_sprite[0][70][24] = 1;dino_sprite[0][70][25] = 1;dino_sprite[0][70][26] = 1;dino_sprite[0][70][27] = 1;dino_sprite[0][70][28] = 1;dino_sprite[0][70][29] = 1;dino_sprite[0][70][30] = 1;dino_sprite[0][70][31] = 1;dino_sprite[0][70][32] = 1;dino_sprite[0][70][33] = 1;dino_sprite[0][70][34] = 1;dino_sprite[0][70][35] = 1;dino_sprite[0][70][36] = 1;dino_sprite[0][70][37] = 1;dino_sprite[0][70][38] = 1;dino_sprite[0][70][39] = 1;dino_sprite[0][70][40] = 1;dino_sprite[0][70][41] = 1;dino_sprite[0][70][42] = 1;dino_sprite[0][70][43] = 1;dino_sprite[0][70][44] = 1;dino_sprite[0][70][45] = 1;dino_sprite[0][70][46] = 1;dino_sprite[0][70][47] = 1;dino_sprite[0][70][48] = 1;dino_sprite[0][70][49] = 1;dino_sprite[0][70][50] = 1;dino_sprite[0][70][51] = 1;dino_sprite[0][70][52] = 1;dino_sprite[0][70][53] = 1;dino_sprite[0][70][54] = 1;dino_sprite[0][70][55] = 1;dino_sprite[0][70][56] = 1;dino_sprite[0][70][57] = 1;dino_sprite[0][70][58] = 1;dino_sprite[0][70][59] = 1;dino_sprite[0][70][60] = 1;dino_sprite[0][70][61] = 1;dino_sprite[0][70][62] = 1;dino_sprite[0][70][63] = 1;dino_sprite[0][70][64] = 1;dino_sprite[0][70][65] = 1;dino_sprite[0][71][0] = 1;dino_sprite[0][71][1] = 1;dino_sprite[0][71][2] = 1;dino_sprite[0][71][3] = 1;dino_sprite[0][71][4] = 1;dino_sprite[0][71][5] = 1;dino_sprite[0][71][6] = 1;dino_sprite[0][71][7] = 1;dino_sprite[0][71][8] = 1;dino_sprite[0][71][9] = 1;dino_sprite[0][71][10] = 1;dino_sprite[0][71][11] = 1;dino_sprite[0][71][12] = 1;dino_sprite[0][71][13] = 1;dino_sprite[0][71][14] = 1;dino_sprite[0][71][15] = 1;dino_sprite[0][71][16] = 1;dino_sprite[0][71][17] = 1;dino_sprite[0][71][18] = 1;dino_sprite[0][71][19] = 1;dino_sprite[0][71][20] = 1;dino_sprite[0][71][21] = 1;dino_sprite[0][71][22] = 1;dino_sprite[0][71][23] = 1;dino_sprite[0][71][24] = 1;dino_sprite[0][71][25] = 1;dino_sprite[0][71][26] = 1;dino_sprite[0][71][27] = 1;dino_sprite[0][71][28] = 1;dino_sprite[0][71][29] = 1;dino_sprite[0][71][30] = 1;dino_sprite[0][71][31] = 1;dino_sprite[0][71][32] = 1;dino_sprite[0][71][33] = 1;dino_sprite[0][71][34] = 1;dino_sprite[0][71][35] = 1;dino_sprite[0][71][36] = 1;dino_sprite[0][71][37] = 1;dino_sprite[0][71][38] = 1;dino_sprite[0][71][39] = 1;dino_sprite[0][71][40] = 1;dino_sprite[0][71][41] = 1;dino_sprite[0][71][43] = 1;dino_sprite[0][71][44] = 1;dino_sprite[0][71][45] = 1;dino_sprite[0][71][46] = 1;dino_sprite[0][71][47] = 1;dino_sprite[0][71][48] = 1;dino_sprite[0][71][49] = 1;dino_sprite[0][72][0] = 1;dino_sprite[0][72][1] = 1;dino_sprite[0][72][2] = 1;dino_sprite[0][72][3] = 1;dino_sprite[0][72][4] = 1;dino_sprite[0][72][5] = 1;dino_sprite[0][72][6] = 1;dino_sprite[0][72][7] = 1;dino_sprite[0][72][8] = 1;dino_sprite[0][72][9] = 1;dino_sprite[0][72][10] = 1;dino_sprite[0][72][11] = 1;dino_sprite[0][72][12] = 1;dino_sprite[0][72][13] = 1;dino_sprite[0][72][14] = 1;dino_sprite[0][72][15] = 1;dino_sprite[0][72][16] = 1;dino_sprite[0][72][17] = 1;dino_sprite[0][72][18] = 1;dino_sprite[0][72][19] = 1;dino_sprite[0][72][20] = 1;dino_sprite[0][72][21] = 1;dino_sprite[0][72][22] = 1;dino_sprite[0][72][23] = 1;dino_sprite[0][72][24] = 1;dino_sprite[0][72][25] = 1;dino_sprite[0][72][26] = 1;dino_sprite[0][72][27] = 1;dino_sprite[0][72][28] = 1;dino_sprite[0][72][29] = 1;dino_sprite[0][72][30] = 1;dino_sprite[0][72][31] = 1;dino_sprite[0][72][32] = 1;dino_sprite[0][72][33] = 1;dino_sprite[0][72][34] = 1;dino_sprite[0][72][35] = 1;dino_sprite[0][72][43] = 1;dino_sprite[0][72][44] = 1;dino_sprite[0][72][45] = 1;dino_sprite[0][72][46] = 1;dino_sprite[0][72][47] = 1;dino_sprite[0][72][48] = 1;dino_sprite[0][72][49] = 1;dino_sprite[0][73][0] = 1;dino_sprite[0][73][1] = 1;dino_sprite[0][73][2] = 1;dino_sprite[0][73][3] = 1;dino_sprite[0][73][4] = 1;dino_sprite[0][73][5] = 1;dino_sprite[0][73][6] = 1;dino_sprite[0][73][7] = 1;dino_sprite[0][73][8] = 1;dino_sprite[0][73][9] = 1;dino_sprite[0][73][10] = 1;dino_sprite[0][73][11] = 1;dino_sprite[0][73][12] = 1;dino_sprite[0][73][13] = 1;dino_sprite[0][73][14] = 1;dino_sprite[0][73][15] = 1;dino_sprite[0][73][16] = 1;dino_sprite[0][73][17] = 1;dino_sprite[0][73][18] = 1;dino_sprite[0][73][19] = 1;dino_sprite[0][73][20] = 1;dino_sprite[0][73][21] = 1;dino_sprite[0][73][22] = 1;dino_sprite[0][73][23] = 1;dino_sprite[0][73][24] = 1;dino_sprite[0][73][25] = 1;dino_sprite[0][73][26] = 1;dino_sprite[0][73][27] = 1;dino_sprite[0][73][28] = 1;dino_sprite[0][73][29] = 1;dino_sprite[0][73][30] = 1;dino_sprite[0][73][31] = 1;dino_sprite[0][73][32] = 1;dino_sprite[0][73][33] = 1;dino_sprite[0][73][34] = 1;dino_sprite[0][73][35] = 1;dino_sprite[0][73][43] = 1;dino_sprite[0][73][44] = 1;dino_sprite[0][73][45] = 1;dino_sprite[0][73][46] = 1;dino_sprite[0][73][47] = 1;dino_sprite[0][73][48] = 1;dino_sprite[0][73][49] = 1;dino_sprite[0][74][0] = 1;dino_sprite[0][74][1] = 1;dino_sprite[0][74][2] = 1;dino_sprite[0][74][3] = 1;dino_sprite[0][74][4] = 1;dino_sprite[0][74][5] = 1;dino_sprite[0][74][6] = 1;dino_sprite[0][74][7] = 1;dino_sprite[0][74][8] = 1;dino_sprite[0][74][9] = 1;dino_sprite[0][74][10] = 1;dino_sprite[0][74][11] = 1;dino_sprite[0][74][12] = 1;dino_sprite[0][74][13] = 1;dino_sprite[0][74][14] = 1;dino_sprite[0][74][15] = 1;dino_sprite[0][74][16] = 1;dino_sprite[0][74][17] = 1;dino_sprite[0][74][18] = 1;dino_sprite[0][74][19] = 1;dino_sprite[0][74][20] = 1;dino_sprite[0][74][21] = 1;dino_sprite[0][74][22] = 1;dino_sprite[0][74][23] = 1;dino_sprite[0][74][24] = 1;dino_sprite[0][74][25] = 1;dino_sprite[0][74][26] = 1;dino_sprite[0][74][27] = 1;dino_sprite[0][74][28] = 1;dino_sprite[0][74][29] = 1;dino_sprite[0][74][30] = 1;dino_sprite[0][74][31] = 1;dino_sprite[0][74][32] = 1;dino_sprite[0][74][33] = 1;dino_sprite[0][74][34] = 1;dino_sprite[0][74][35] = 1;dino_sprite[0][74][43] = 1;dino_sprite[0][74][44] = 1;dino_sprite[0][74][45] = 1;dino_sprite[0][74][46] = 1;dino_sprite[0][74][47] = 1;dino_sprite[0][74][48] = 1;dino_sprite[0][74][49] = 1;dino_sprite[0][75][0] = 1;dino_sprite[0][75][1] = 1;dino_sprite[0][75][2] = 1;dino_sprite[0][75][3] = 1;dino_sprite[0][75][4] = 1;dino_sprite[0][75][5] = 1;dino_sprite[0][75][6] = 1;dino_sprite[0][75][7] = 1;dino_sprite[0][75][8] = 1;dino_sprite[0][75][9] = 1;dino_sprite[0][75][10] = 1;dino_sprite[0][75][11] = 1;dino_sprite[0][75][12] = 1;dino_sprite[0][75][13] = 1;dino_sprite[0][75][14] = 1;dino_sprite[0][75][15] = 1;dino_sprite[0][75][16] = 1;dino_sprite[0][75][17] = 1;dino_sprite[0][75][18] = 1;dino_sprite[0][75][19] = 1;dino_sprite[0][75][20] = 1;dino_sprite[0][75][21] = 1;dino_sprite[0][75][22] = 1;dino_sprite[0][75][23] = 1;dino_sprite[0][75][24] = 1;dino_sprite[0][75][25] = 1;dino_sprite[0][75][26] = 1;dino_sprite[0][75][27] = 1;dino_sprite[0][75][28] = 1;dino_sprite[0][75][29] = 1;dino_sprite[0][75][30] = 1;dino_sprite[0][75][31] = 1;dino_sprite[0][75][32] = 1;dino_sprite[0][75][33] = 1;dino_sprite[0][75][34] = 1;dino_sprite[0][75][35] = 1;dino_sprite[0][75][43] = 1;dino_sprite[0][75][44] = 1;dino_sprite[0][75][45] = 1;dino_sprite[0][75][46] = 1;dino_sprite[0][75][47] = 1;dino_sprite[0][75][48] = 1;dino_sprite[0][75][49] = 1;dino_sprite[0][75][50] = 1;dino_sprite[0][75][51] = 1;dino_sprite[0][75][52] = 1;dino_sprite[0][75][53] = 1;dino_sprite[0][75][54] = 1;dino_sprite[0][76][0] = 1;dino_sprite[0][76][1] = 1;dino_sprite[0][76][2] = 1;dino_sprite[0][76][3] = 1;dino_sprite[0][76][4] = 1;dino_sprite[0][76][5] = 1;dino_sprite[0][76][6] = 1;dino_sprite[0][76][7] = 1;dino_sprite[0][76][8] = 1;dino_sprite[0][76][9] = 1;dino_sprite[0][76][10] = 1;dino_sprite[0][76][11] = 1;dino_sprite[0][76][12] = 1;dino_sprite[0][76][13] = 1;dino_sprite[0][76][14] = 1;dino_sprite[0][76][15] = 1;dino_sprite[0][76][16] = 1;dino_sprite[0][76][17] = 1;dino_sprite[0][76][18] = 1;dino_sprite[0][76][19] = 1;dino_sprite[0][76][20] = 1;dino_sprite[0][76][21] = 1;dino_sprite[0][76][22] = 1;dino_sprite[0][76][23] = 1;dino_sprite[0][76][24] = 1;dino_sprite[0][76][25] = 1;dino_sprite[0][76][26] = 1;dino_sprite[0][76][27] = 1;dino_sprite[0][76][28] = 1;dino_sprite[0][76][29] = 1;dino_sprite[0][76][30] = 1;dino_sprite[0][76][31] = 1;dino_sprite[0][76][32] = 1;dino_sprite[0][76][33] = 1;dino_sprite[0][76][34] = 1;dino_sprite[0][76][35] = 1;dino_sprite[0][76][43] = 1;dino_sprite[0][76][44] = 1;dino_sprite[0][76][45] = 1;dino_sprite[0][76][46] = 1;dino_sprite[0][76][47] = 1;dino_sprite[0][76][48] = 1;dino_sprite[0][76][49] = 1;dino_sprite[0][76][50] = 1;dino_sprite[0][76][51] = 1;dino_sprite[0][76][52] = 1;dino_sprite[0][76][53] = 1;dino_sprite[0][76][54] = 1;dino_sprite[0][77][0] = 1;dino_sprite[0][77][1] = 1;dino_sprite[0][77][2] = 1;dino_sprite[0][77][3] = 1;dino_sprite[0][77][4] = 1;dino_sprite[0][77][5] = 1;dino_sprite[0][77][6] = 1;dino_sprite[0][77][7] = 1;dino_sprite[0][77][8] = 1;dino_sprite[0][77][9] = 1;dino_sprite[0][77][10] = 1;dino_sprite[0][77][11] = 1;dino_sprite[0][77][12] = 1;dino_sprite[0][77][13] = 1;dino_sprite[0][77][14] = 1;dino_sprite[0][77][15] = 1;dino_sprite[0][77][16] = 1;dino_sprite[0][77][17] = 1;dino_sprite[0][77][18] = 1;dino_sprite[0][77][19] = 1;dino_sprite[0][77][20] = 1;dino_sprite[0][77][21] = 1;dino_sprite[0][77][22] = 1;dino_sprite[0][77][23] = 1;dino_sprite[0][77][24] = 1;dino_sprite[0][77][25] = 1;dino_sprite[0][77][29] = 1;dino_sprite[0][77][30] = 1;dino_sprite[0][77][31] = 1;dino_sprite[0][77][32] = 1;dino_sprite[0][77][33] = 1;dino_sprite[0][77][34] = 1;dino_sprite[0][77][35] = 1;dino_sprite[0][77][43] = 1;dino_sprite[0][77][44] = 1;dino_sprite[0][77][45] = 1;dino_sprite[0][77][46] = 1;dino_sprite[0][77][47] = 1;dino_sprite[0][77][48] = 1;dino_sprite[0][77][49] = 1;dino_sprite[0][77][50] = 1;dino_sprite[0][77][51] = 1;dino_sprite[0][77][52] = 1;dino_sprite[0][77][53] = 1;dino_sprite[0][77][54] = 1;dino_sprite[0][78][0] = 1;dino_sprite[0][78][1] = 1;dino_sprite[0][78][2] = 1;dino_sprite[0][78][3] = 1;dino_sprite[0][78][4] = 1;dino_sprite[0][78][5] = 1;dino_sprite[0][78][6] = 1;dino_sprite[0][78][7] = 1;dino_sprite[0][78][8] = 1;dino_sprite[0][78][9] = 1;dino_sprite[0][78][10] = 1;dino_sprite[0][78][11] = 1;dino_sprite[0][78][12] = 1;dino_sprite[0][78][13] = 1;dino_sprite[0][78][14] = 1;dino_sprite[0][78][15] = 1;dino_sprite[0][78][16] = 1;dino_sprite[0][78][17] = 1;dino_sprite[0][78][18] = 1;dino_sprite[0][78][19] = 1;dino_sprite[0][78][20] = 1;dino_sprite[0][78][21] = 1;dino_sprite[0][78][22] = 1;dino_sprite[0][78][23] = 1;dino_sprite[0][78][24] = 1;dino_sprite[0][78][25] = 1;dino_sprite[0][78][29] = 1;dino_sprite[0][78][30] = 1;dino_sprite[0][78][31] = 1;dino_sprite[0][78][32] = 1;dino_sprite[0][78][33] = 1;dino_sprite[0][78][34] = 1;dino_sprite[0][78][35] = 1;dino_sprite[0][78][43] = 1;dino_sprite[0][78][44] = 1;dino_sprite[0][78][45] = 1;dino_sprite[0][78][46] = 1;dino_sprite[0][78][47] = 1;dino_sprite[0][78][48] = 1;dino_sprite[0][78][49] = 1;dino_sprite[0][78][50] = 1;dino_sprite[0][78][51] = 1;dino_sprite[0][78][52] = 1;dino_sprite[0][78][53] = 1;dino_sprite[0][78][54] = 1;dino_sprite[0][79][0] = 1;dino_sprite[0][79][1] = 1;dino_sprite[0][79][2] = 1;dino_sprite[0][79][3] = 1;dino_sprite[0][79][4] = 1;dino_sprite[0][79][5] = 1;dino_sprite[0][79][6] = 1;dino_sprite[0][79][7] = 1;dino_sprite[0][79][8] = 1;dino_sprite[0][79][9] = 1;dino_sprite[0][79][10] = 1;dino_sprite[0][79][11] = 1;dino_sprite[0][79][12] = 1;dino_sprite[0][79][13] = 1;dino_sprite[0][79][14] = 1;dino_sprite[0][79][15] = 1;dino_sprite[0][79][16] = 1;dino_sprite[0][79][17] = 1;dino_sprite[0][79][18] = 1;dino_sprite[0][79][19] = 1;dino_sprite[0][79][20] = 1;dino_sprite[0][79][21] = 1;dino_sprite[0][79][22] = 1;dino_sprite[0][79][23] = 1;dino_sprite[0][79][24] = 1;dino_sprite[0][79][25] = 1;dino_sprite[0][79][29] = 1;dino_sprite[0][79][30] = 1;dino_sprite[0][79][31] = 1;dino_sprite[0][79][32] = 1;dino_sprite[0][79][33] = 1;dino_sprite[0][79][34] = 1;dino_sprite[0][79][35] = 1;dino_sprite[0][79][43] = 1;dino_sprite[0][79][44] = 1;dino_sprite[0][79][45] = 1;dino_sprite[0][79][46] = 1;dino_sprite[0][79][47] = 1;dino_sprite[0][79][48] = 1;dino_sprite[0][79][49] = 1;dino_sprite[0][79][50] = 1;dino_sprite[0][79][51] = 1;dino_sprite[0][79][52] = 1;dino_sprite[0][79][53] = 1;dino_sprite[0][79][54] = 1;dino_sprite[0][80][0] = 1;dino_sprite[0][80][1] = 1;dino_sprite[0][80][2] = 1;dino_sprite[0][80][3] = 1;dino_sprite[0][80][4] = 1;dino_sprite[0][80][5] = 1;dino_sprite[0][80][6] = 1;dino_sprite[0][80][7] = 1;dino_sprite[0][80][8] = 1;dino_sprite[0][80][9] = 1;dino_sprite[0][80][10] = 1;dino_sprite[0][80][11] = 1;dino_sprite[0][80][12] = 1;dino_sprite[0][80][13] = 1;dino_sprite[0][80][14] = 1;dino_sprite[0][80][15] = 1;dino_sprite[0][80][16] = 1;dino_sprite[0][80][17] = 1;dino_sprite[0][80][18] = 1;dino_sprite[0][80][19] = 1;dino_sprite[0][80][20] = 1;dino_sprite[0][80][21] = 1;dino_sprite[0][80][22] = 1;dino_sprite[0][80][23] = 1;dino_sprite[0][80][24] = 1;dino_sprite[0][80][25] = 1;dino_sprite[0][80][29] = 1;dino_sprite[0][80][30] = 1;dino_sprite[0][80][31] = 1;dino_sprite[0][80][32] = 1;dino_sprite[0][80][33] = 1;dino_sprite[0][80][34] = 1;dino_sprite[0][80][35] = 1;dino_sprite[0][80][43] = 1;dino_sprite[0][80][44] = 1;dino_sprite[0][80][45] = 1;dino_sprite[0][80][46] = 1;dino_sprite[0][80][47] = 1;dino_sprite[0][80][48] = 1;dino_sprite[0][80][49] = 1;dino_sprite[0][80][50] = 1;dino_sprite[0][80][51] = 1;dino_sprite[0][80][52] = 1;dino_sprite[0][80][53] = 1;dino_sprite[0][80][54] = 1;dino_sprite[0][81][0] = 1;dino_sprite[0][81][1] = 1;dino_sprite[0][81][2] = 1;dino_sprite[0][81][3] = 1;dino_sprite[0][81][4] = 1;dino_sprite[0][81][5] = 1;dino_sprite[0][81][6] = 1;dino_sprite[0][81][7] = 1;dino_sprite[0][81][8] = 1;dino_sprite[0][81][9] = 1;dino_sprite[0][81][10] = 1;dino_sprite[0][81][11] = 1;dino_sprite[0][81][12] = 1;dino_sprite[0][81][13] = 1;dino_sprite[0][81][14] = 1;dino_sprite[0][81][15] = 1;dino_sprite[0][81][16] = 1;dino_sprite[0][81][17] = 1;dino_sprite[0][81][18] = 1;dino_sprite[0][81][19] = 1;dino_sprite[0][81][20] = 1;dino_sprite[0][81][21] = 1;dino_sprite[0][81][22] = 1;dino_sprite[0][81][23] = 1;dino_sprite[0][81][24] = 1;dino_sprite[0][81][25] = 1;dino_sprite[0][81][29] = 1;dino_sprite[0][81][30] = 1;dino_sprite[0][81][31] = 1;dino_sprite[0][81][32] = 1;dino_sprite[0][81][33] = 1;dino_sprite[0][81][34] = 1;dino_sprite[0][81][35] = 1;dino_sprite[0][81][43] = 1;dino_sprite[0][81][44] = 1;dino_sprite[0][81][45] = 1;dino_sprite[0][81][46] = 1;dino_sprite[0][81][47] = 1;dino_sprite[0][81][48] = 1;dino_sprite[0][81][49] = 1;dino_sprite[0][81][50] = 1;dino_sprite[0][81][51] = 1;dino_sprite[0][81][52] = 1;dino_sprite[0][81][53] = 1;dino_sprite[0][81][54] = 1;dino_sprite[0][82][0] = 1;dino_sprite[0][82][1] = 1;dino_sprite[0][82][2] = 1;dino_sprite[0][82][3] = 1;dino_sprite[0][82][4] = 1;dino_sprite[0][82][5] = 1;dino_sprite[0][82][6] = 1;dino_sprite[0][82][7] = 1;dino_sprite[0][82][8] = 1;dino_sprite[0][82][9] = 1;dino_sprite[0][82][10] = 1;dino_sprite[0][82][11] = 1;dino_sprite[0][82][12] = 1;dino_sprite[0][82][13] = 1;dino_sprite[0][82][14] = 1;dino_sprite[0][82][15] = 1;dino_sprite[0][82][16] = 1;dino_sprite[0][82][17] = 1;dino_sprite[0][82][18] = 1;dino_sprite[0][82][19] = 1;dino_sprite[0][82][20] = 1;dino_sprite[0][82][21] = 1;dino_sprite[0][82][22] = 1;dino_sprite[0][82][23] = 1;dino_sprite[0][82][24] = 1;dino_sprite[0][82][25] = 1;dino_sprite[0][82][29] = 1;dino_sprite[0][82][30] = 1;dino_sprite[0][82][31] = 1;dino_sprite[0][82][32] = 1;dino_sprite[0][82][33] = 1;dino_sprite[0][82][34] = 1;dino_sprite[0][82][35] = 1;dino_sprite[0][83][0] = 1;dino_sprite[0][83][1] = 1;dino_sprite[0][83][2] = 1;dino_sprite[0][83][3] = 1;dino_sprite[0][83][4] = 1;dino_sprite[0][83][5] = 1;dino_sprite[0][83][6] = 1;dino_sprite[0][83][7] = 1;dino_sprite[0][83][8] = 1;dino_sprite[0][83][9] = 1;dino_sprite[0][83][10] = 1;dino_sprite[0][83][11] = 1;dino_sprite[0][83][12] = 1;dino_sprite[0][83][13] = 1;dino_sprite[0][83][14] = 1;dino_sprite[0][83][15] = 1;dino_sprite[0][83][16] = 1;dino_sprite[0][83][17] = 1;dino_sprite[0][83][18] = 1;dino_sprite[0][83][19] = 1;dino_sprite[0][83][20] = 1;dino_sprite[0][83][21] = 1;dino_sprite[0][83][22] = 1;dino_sprite[0][83][23] = 1;dino_sprite[0][83][24] = 1;dino_sprite[0][83][25] = 1;dino_sprite[0][83][29] = 1;dino_sprite[0][83][30] = 1;dino_sprite[0][83][31] = 1;dino_sprite[0][83][32] = 1;dino_sprite[0][83][33] = 1;dino_sprite[0][83][34] = 1;dino_sprite[0][83][35] = 1;dino_sprite[0][84][0] = 1;dino_sprite[0][84][1] = 1;dino_sprite[0][84][2] = 1;dino_sprite[0][84][3] = 1;dino_sprite[0][84][4] = 1;dino_sprite[0][84][5] = 1;dino_sprite[0][84][6] = 1;dino_sprite[0][84][7] = 1;dino_sprite[0][84][8] = 1;dino_sprite[0][84][9] = 1;dino_sprite[0][84][10] = 1;dino_sprite[0][84][11] = 1;dino_sprite[0][84][12] = 1;dino_sprite[0][84][13] = 1;dino_sprite[0][84][14] = 1;dino_sprite[0][84][15] = 1;dino_sprite[0][84][16] = 1;dino_sprite[0][84][17] = 1;dino_sprite[0][84][18] = 1;dino_sprite[0][84][19] = 1;dino_sprite[0][84][20] = 1;dino_sprite[0][84][21] = 1;dino_sprite[0][84][22] = 1;dino_sprite[0][84][23] = 1;dino_sprite[0][84][24] = 1;dino_sprite[0][84][25] = 1;dino_sprite[0][84][29] = 1;dino_sprite[0][84][30] = 1;dino_sprite[0][84][31] = 1;dino_sprite[0][84][32] = 1;dino_sprite[0][84][33] = 1;dino_sprite[0][84][34] = 1;dino_sprite[0][84][35] = 1;dino_sprite[0][85][0] = 1;dino_sprite[0][85][1] = 1;dino_sprite[0][85][2] = 1;dino_sprite[0][85][3] = 1;dino_sprite[0][85][4] = 1;dino_sprite[0][85][5] = 1;dino_sprite[0][85][6] = 1;dino_sprite[0][85][7] = 1;dino_sprite[0][85][8] = 1;dino_sprite[0][85][9] = 1;dino_sprite[0][85][10] = 1;dino_sprite[0][85][11] = 1;dino_sprite[0][85][12] = 1;dino_sprite[0][85][13] = 1;dino_sprite[0][85][14] = 1;dino_sprite[0][85][15] = 1;dino_sprite[0][85][16] = 1;dino_sprite[0][85][17] = 1;dino_sprite[0][85][18] = 1;dino_sprite[0][85][19] = 1;dino_sprite[0][85][20] = 1;dino_sprite[0][85][21] = 1;dino_sprite[0][85][22] = 1;dino_sprite[0][85][23] = 1;dino_sprite[0][85][24] = 1;dino_sprite[0][85][25] = 1;dino_sprite[0][85][29] = 1;dino_sprite[0][85][30] = 1;dino_sprite[0][85][31] = 1;dino_sprite[0][85][32] = 1;dino_sprite[0][85][33] = 1;dino_sprite[0][85][34] = 1;dino_sprite[0][85][35] = 1;dino_sprite[0][86][0] = 1;dino_sprite[0][86][1] = 1;dino_sprite[0][86][2] = 1;dino_sprite[0][86][3] = 1;dino_sprite[0][86][4] = 1;dino_sprite[0][86][5] = 1;dino_sprite[0][86][6] = 1;dino_sprite[0][86][7] = 1;dino_sprite[0][86][8] = 1;dino_sprite[0][86][9] = 1;dino_sprite[0][86][10] = 1;dino_sprite[0][86][11] = 1;dino_sprite[0][86][12] = 1;dino_sprite[0][86][13] = 1;dino_sprite[0][86][14] = 1;dino_sprite[0][86][15] = 1;dino_sprite[0][86][16] = 1;dino_sprite[0][86][17] = 1;dino_sprite[0][86][18] = 1;dino_sprite[0][86][19] = 1;dino_sprite[0][86][20] = 1;dino_sprite[0][86][21] = 1;dino_sprite[0][86][22] = 1;dino_sprite[0][86][23] = 1;dino_sprite[0][86][24] = 1;dino_sprite[0][86][25] = 1;dino_sprite[0][86][29] = 1;dino_sprite[0][86][30] = 1;dino_sprite[0][86][31] = 1;dino_sprite[0][86][32] = 1;dino_sprite[0][86][33] = 1;dino_sprite[0][86][34] = 1;dino_sprite[0][86][35] = 1;dino_sprite[0][87][0] = 1;dino_sprite[0][87][1] = 1;dino_sprite[0][87][2] = 1;dino_sprite[0][87][3] = 1;dino_sprite[0][87][4] = 1;dino_sprite[0][87][5] = 1;dino_sprite[0][87][6] = 1;dino_sprite[0][87][7] = 1;dino_sprite[0][87][8] = 1;dino_sprite[0][87][9] = 1;dino_sprite[0][87][10] = 1;dino_sprite[0][87][11] = 1;dino_sprite[0][87][12] = 1;dino_sprite[0][87][13] = 1;dino_sprite[0][87][14] = 1;dino_sprite[0][87][15] = 1;dino_sprite[0][87][16] = 1;dino_sprite[0][87][17] = 1;dino_sprite[0][87][18] = 1;dino_sprite[0][87][19] = 1;dino_sprite[0][87][20] = 1;dino_sprite[0][87][21] = 1;dino_sprite[0][87][22] = 1;dino_sprite[0][87][23] = 1;dino_sprite[0][87][24] = 1;dino_sprite[0][87][25] = 1;dino_sprite[0][87][29] = 1;dino_sprite[0][87][30] = 1;dino_sprite[0][87][31] = 1;dino_sprite[0][87][32] = 1;dino_sprite[0][87][33] = 1;dino_sprite[0][87][34] = 1;dino_sprite[0][87][35] = 1;dino_sprite[0][88][0] = 1;dino_sprite[0][88][1] = 1;dino_sprite[0][88][2] = 1;dino_sprite[0][88][3] = 1;dino_sprite[0][88][4] = 1;dino_sprite[0][88][5] = 1;dino_sprite[0][88][6] = 1;dino_sprite[0][88][7] = 1;dino_sprite[0][88][8] = 1;dino_sprite[0][88][9] = 1;dino_sprite[0][88][10] = 1;dino_sprite[0][88][11] = 1;dino_sprite[0][88][12] = 1;dino_sprite[0][88][13] = 1;dino_sprite[0][88][14] = 1;dino_sprite[0][88][15] = 1;dino_sprite[0][88][16] = 1;dino_sprite[0][88][17] = 1;dino_sprite[0][88][18] = 1;dino_sprite[0][88][19] = 1;dino_sprite[0][88][20] = 1;dino_sprite[0][88][21] = 1;dino_sprite[0][88][22] = 1;dino_sprite[0][88][23] = 1;dino_sprite[0][88][24] = 1;dino_sprite[0][88][25] = 1;dino_sprite[0][88][29] = 1;dino_sprite[0][88][30] = 1;dino_sprite[0][88][31] = 1;dino_sprite[0][88][32] = 1;dino_sprite[0][88][33] = 1;dino_sprite[0][88][34] = 1;dino_sprite[0][88][35] = 1;dino_sprite[0][89][0] = 1;dino_sprite[0][89][1] = 1;dino_sprite[0][89][2] = 1;dino_sprite[0][89][3] = 1;dino_sprite[0][89][4] = 1;dino_sprite[0][89][5] = 1;dino_sprite[0][89][6] = 1;dino_sprite[0][89][7] = 1;dino_sprite[0][89][8] = 1;dino_sprite[0][89][9] = 1;dino_sprite[0][89][10] = 1;dino_sprite[0][89][11] = 1;dino_sprite[0][89][12] = 1;dino_sprite[0][89][13] = 1;dino_sprite[0][89][14] = 1;dino_sprite[0][89][15] = 1;dino_sprite[0][89][16] = 1;dino_sprite[0][89][17] = 1;dino_sprite[0][89][18] = 1;dino_sprite[0][89][19] = 1;dino_sprite[0][89][20] = 1;dino_sprite[0][89][21] = 1;dino_sprite[0][89][22] = 1;dino_sprite[0][89][23] = 1;dino_sprite[0][89][24] = 1;dino_sprite[0][89][25] = 1;dino_sprite[0][89][29] = 1;dino_sprite[0][89][30] = 1;dino_sprite[0][89][31] = 1;dino_sprite[0][89][32] = 1;dino_sprite[0][89][33] = 1;dino_sprite[0][89][34] = 1;dino_sprite[0][89][35] = 1;dino_sprite[0][90][0] = 1;dino_sprite[0][90][1] = 1;dino_sprite[0][90][2] = 1;dino_sprite[0][90][3] = 1;dino_sprite[0][90][4] = 1;dino_sprite[0][90][5] = 1;dino_sprite[0][90][6] = 1;dino_sprite[0][90][7] = 1;dino_sprite[0][90][8] = 1;dino_sprite[0][90][9] = 1;dino_sprite[0][90][10] = 1;dino_sprite[0][90][11] = 1;dino_sprite[0][90][12] = 1;dino_sprite[0][90][13] = 1;dino_sprite[0][90][14] = 1;dino_sprite[0][90][15] = 1;dino_sprite[0][90][16] = 1;dino_sprite[0][90][17] = 1;dino_sprite[0][90][18] = 1;dino_sprite[0][90][19] = 1;dino_sprite[0][90][20] = 1;dino_sprite[0][90][21] = 1;dino_sprite[0][90][22] = 1;dino_sprite[0][90][23] = 1;dino_sprite[0][90][24] = 1;dino_sprite[0][90][25] = 1;dino_sprite[0][90][29] = 1;dino_sprite[0][90][30] = 1;dino_sprite[0][90][31] = 1;dino_sprite[0][90][32] = 1;dino_sprite[0][90][33] = 1;dino_sprite[0][90][34] = 1;dino_sprite[0][90][35] = 1;dino_sprite[0][91][0] = 1;dino_sprite[0][91][1] = 1;dino_sprite[0][91][2] = 1;dino_sprite[0][91][3] = 1;dino_sprite[0][91][4] = 1;dino_sprite[0][91][5] = 1;dino_sprite[0][91][6] = 1;dino_sprite[0][91][7] = 1;dino_sprite[0][91][8] = 1;dino_sprite[0][91][9] = 1;dino_sprite[0][91][10] = 1;dino_sprite[0][91][11] = 1;dino_sprite[0][91][12] = 1;dino_sprite[0][91][13] = 1;dino_sprite[0][91][14] = 1;dino_sprite[0][91][15] = 1;dino_sprite[0][91][16] = 1;dino_sprite[0][91][17] = 1;dino_sprite[0][91][18] = 1;dino_sprite[0][91][19] = 1;dino_sprite[0][91][20] = 1;dino_sprite[0][91][21] = 1;dino_sprite[0][91][22] = 1;dino_sprite[0][91][23] = 1;dino_sprite[0][91][24] = 1;dino_sprite[0][91][25] = 1;dino_sprite[0][91][30] = 1;dino_sprite[0][91][31] = 1;dino_sprite[0][91][32] = 1;dino_sprite[0][91][33] = 1;dino_sprite[0][92][0] = 1;dino_sprite[0][92][1] = 1;dino_sprite[0][92][2] = 1;dino_sprite[0][92][3] = 1;dino_sprite[0][92][4] = 1;dino_sprite[0][92][5] = 1;dino_sprite[0][92][6] = 1;dino_sprite[0][92][7] = 1;dino_sprite[0][92][8] = 1;dino_sprite[0][92][9] = 1;dino_sprite[0][92][10] = 1;dino_sprite[0][92][11] = 1;dino_sprite[0][92][12] = 1;dino_sprite[0][92][13] = 1;dino_sprite[0][92][14] = 1;dino_sprite[0][92][15] = 1;dino_sprite[0][92][16] = 1;dino_sprite[0][92][17] = 1;dino_sprite[0][92][18] = 1;dino_sprite[0][92][19] = 1;dino_sprite[0][92][20] = 1;dino_sprite[0][92][21] = 1;dino_sprite[0][92][22] = 1;dino_sprite[0][92][23] = 1;dino_sprite[0][92][24] = 1;dino_sprite[0][92][25] = 1;dino_sprite[0][93][0] = 1;dino_sprite[0][93][1] = 1;dino_sprite[0][93][2] = 1;dino_sprite[0][93][3] = 1;dino_sprite[0][93][4] = 1;dino_sprite[0][93][5] = 1;dino_sprite[0][93][6] = 1;dino_sprite[0][93][7] = 1;dino_sprite[0][93][8] = 1;dino_sprite[0][93][9] = 1;dino_sprite[0][93][10] = 1;dino_sprite[0][93][11] = 1;dino_sprite[0][93][12] = 1;dino_sprite[0][93][13] = 1;dino_sprite[0][93][14] = 1;dino_sprite[0][93][15] = 1;dino_sprite[0][93][16] = 1;dino_sprite[0][93][17] = 1;dino_sprite[0][93][18] = 1;dino_sprite[0][93][19] = 1;dino_sprite[0][93][20] = 1;dino_sprite[0][93][21] = 1;dino_sprite[0][93][22] = 1;dino_sprite[0][93][23] = 1;dino_sprite[0][93][24] = 1;dino_sprite[0][93][25] = 1;dino_sprite[0][94][0] = 1;dino_sprite[0][94][1] = 1;dino_sprite[0][94][2] = 1;dino_sprite[0][94][3] = 1;dino_sprite[0][94][4] = 1;dino_sprite[0][94][5] = 1;dino_sprite[0][94][6] = 1;dino_sprite[0][94][7] = 1;dino_sprite[0][94][8] = 1;dino_sprite[0][94][9] = 1;dino_sprite[0][94][10] = 1;dino_sprite[0][94][11] = 1;dino_sprite[0][94][12] = 1;dino_sprite[0][94][13] = 1;dino_sprite[0][94][14] = 1;dino_sprite[0][94][15] = 1;dino_sprite[0][94][16] = 1;dino_sprite[0][94][17] = 1;dino_sprite[0][94][18] = 1;dino_sprite[0][94][19] = 1;dino_sprite[0][94][20] = 1;dino_sprite[0][94][21] = 1;dino_sprite[0][94][22] = 1;dino_sprite[0][94][23] = 1;dino_sprite[0][94][24] = 1;dino_sprite[0][94][25] = 1;dino_sprite[0][95][0] = 1;dino_sprite[0][95][1] = 1;dino_sprite[0][95][2] = 1;dino_sprite[0][95][3] = 1;dino_sprite[0][95][4] = 1;dino_sprite[0][95][5] = 1;dino_sprite[0][95][6] = 1;dino_sprite[0][95][7] = 1;dino_sprite[0][95][8] = 1;dino_sprite[0][95][9] = 1;dino_sprite[0][95][10] = 1;dino_sprite[0][95][11] = 1;dino_sprite[0][95][12] = 1;dino_sprite[0][95][13] = 1;dino_sprite[0][95][14] = 1;dino_sprite[0][95][15] = 1;dino_sprite[0][95][16] = 1;dino_sprite[0][95][17] = 1;dino_sprite[0][95][18] = 1;dino_sprite[0][95][19] = 1;dino_sprite[0][95][20] = 1;dino_sprite[0][95][21] = 1;dino_sprite[0][95][22] = 1;dino_sprite[0][95][23] = 1;dino_sprite[0][95][24] = 1;dino_sprite[0][95][25] = 1;dino_sprite[0][96][3] = 1;dino_sprite[0][96][4] = 1;dino_sprite[0][96][5] = 1;dino_sprite[0][96][6] = 1;dino_sprite[0][96][7] = 1;dino_sprite[0][96][8] = 1;dino_sprite[0][96][9] = 1;dino_sprite[0][96][10] = 1;dino_sprite[0][96][11] = 1;dino_sprite[0][96][12] = 1;dino_sprite[0][96][13] = 1;dino_sprite[0][96][14] = 1;dino_sprite[0][96][15] = 1;dino_sprite[0][96][16] = 1;dino_sprite[0][96][17] = 1;dino_sprite[0][96][18] = 1;dino_sprite[0][96][19] = 1;dino_sprite[0][96][20] = 1;dino_sprite[0][96][21] = 1;dino_sprite[0][96][22] = 1;dino_sprite[0][96][23] = 1;dino_sprite[0][96][24] = 1;dino_sprite[0][96][25] = 1;dino_sprite[0][97][3] = 1;dino_sprite[0][97][4] = 1;dino_sprite[0][97][5] = 1;dino_sprite[0][97][6] = 1;dino_sprite[0][97][7] = 1;dino_sprite[0][97][8] = 1;dino_sprite[0][97][9] = 1;dino_sprite[0][97][10] = 1;dino_sprite[0][97][11] = 1;dino_sprite[0][97][12] = 1;dino_sprite[0][97][13] = 1;dino_sprite[0][97][14] = 1;dino_sprite[0][97][15] = 1;dino_sprite[0][97][16] = 1;dino_sprite[0][97][17] = 1;dino_sprite[0][97][18] = 1;dino_sprite[0][97][19] = 1;dino_sprite[0][97][20] = 1;dino_sprite[0][97][21] = 1;dino_sprite[0][97][22] = 1;dino_sprite[0][97][23] = 1;dino_sprite[0][97][24] = 1;dino_sprite[0][97][25] = 1;dino_sprite[0][98][3] = 1;dino_sprite[0][98][4] = 1;dino_sprite[0][98][5] = 1;dino_sprite[0][98][6] = 1;dino_sprite[0][98][7] = 1;dino_sprite[0][98][8] = 1;dino_sprite[0][98][9] = 1;dino_sprite[0][98][10] = 1;dino_sprite[0][98][11] = 1;dino_sprite[0][98][12] = 1;dino_sprite[0][98][13] = 1;dino_sprite[0][98][14] = 1;dino_sprite[0][98][15] = 1;dino_sprite[0][98][16] = 1;dino_sprite[0][98][17] = 1;dino_sprite[0][98][18] = 1;dino_sprite[0][98][19] = 1;dino_sprite[0][98][20] = 1;dino_sprite[0][98][21] = 1;dino_sprite[0][98][22] = 1;dino_sprite[0][98][23] = 1;dino_sprite[0][98][24] = 1;dino_sprite[0][98][25] = 1;
	dino_sprite[1][2][35] = 1;dino_sprite[1][2][36] = 1;dino_sprite[1][2][37] = 1;dino_sprite[1][2][38] = 1;dino_sprite[1][2][39] = 1;dino_sprite[1][2][40] = 1;dino_sprite[1][2][41] = 1;dino_sprite[1][2][42] = 1;dino_sprite[1][2][43] = 1;dino_sprite[1][2][44] = 1;dino_sprite[1][2][45] = 1;dino_sprite[1][2][46] = 1;dino_sprite[1][2][47] = 1;dino_sprite[1][2][48] = 1;dino_sprite[1][2][49] = 1;dino_sprite[1][2][50] = 1;dino_sprite[1][2][51] = 1;dino_sprite[1][2][52] = 1;dino_sprite[1][2][53] = 1;dino_sprite[1][2][54] = 1;dino_sprite[1][2][55] = 1;dino_sprite[1][2][56] = 1;dino_sprite[1][2][57] = 1;dino_sprite[1][2][58] = 1;dino_sprite[1][2][59] = 1;dino_sprite[1][2][60] = 1;dino_sprite[1][2][61] = 1;dino_sprite[1][2][62] = 1;dino_sprite[1][3][35] = 1;dino_sprite[1][3][36] = 1;dino_sprite[1][3][37] = 1;dino_sprite[1][3][38] = 1;dino_sprite[1][3][39] = 1;dino_sprite[1][3][40] = 1;dino_sprite[1][3][41] = 1;dino_sprite[1][3][42] = 1;dino_sprite[1][3][43] = 1;dino_sprite[1][3][44] = 1;dino_sprite[1][3][45] = 1;dino_sprite[1][3][46] = 1;dino_sprite[1][3][47] = 1;dino_sprite[1][3][48] = 1;dino_sprite[1][3][49] = 1;dino_sprite[1][3][50] = 1;dino_sprite[1][3][51] = 1;dino_sprite[1][3][52] = 1;dino_sprite[1][3][53] = 1;dino_sprite[1][3][54] = 1;dino_sprite[1][3][55] = 1;dino_sprite[1][3][56] = 1;dino_sprite[1][3][57] = 1;dino_sprite[1][3][58] = 1;dino_sprite[1][3][59] = 1;dino_sprite[1][3][60] = 1;dino_sprite[1][3][61] = 1;dino_sprite[1][3][62] = 1;dino_sprite[1][4][35] = 1;dino_sprite[1][4][36] = 1;dino_sprite[1][4][37] = 1;dino_sprite[1][4][38] = 1;dino_sprite[1][4][39] = 1;dino_sprite[1][4][40] = 1;dino_sprite[1][4][41] = 1;dino_sprite[1][4][42] = 1;dino_sprite[1][4][43] = 1;dino_sprite[1][4][44] = 1;dino_sprite[1][4][45] = 1;dino_sprite[1][4][46] = 1;dino_sprite[1][4][47] = 1;dino_sprite[1][4][48] = 1;dino_sprite[1][4][49] = 1;dino_sprite[1][4][50] = 1;dino_sprite[1][4][51] = 1;dino_sprite[1][4][52] = 1;dino_sprite[1][4][53] = 1;dino_sprite[1][4][54] = 1;dino_sprite[1][4][55] = 1;dino_sprite[1][4][56] = 1;dino_sprite[1][4][57] = 1;dino_sprite[1][4][58] = 1;dino_sprite[1][4][59] = 1;dino_sprite[1][4][60] = 1;dino_sprite[1][4][61] = 1;dino_sprite[1][4][62] = 1;dino_sprite[1][5][35] = 1;dino_sprite[1][5][36] = 1;dino_sprite[1][5][37] = 1;dino_sprite[1][5][38] = 1;dino_sprite[1][5][39] = 1;dino_sprite[1][5][40] = 1;dino_sprite[1][5][41] = 1;dino_sprite[1][5][42] = 1;dino_sprite[1][5][43] = 1;dino_sprite[1][5][44] = 1;dino_sprite[1][5][45] = 1;dino_sprite[1][5][46] = 1;dino_sprite[1][5][47] = 1;dino_sprite[1][5][48] = 1;dino_sprite[1][5][49] = 1;dino_sprite[1][5][50] = 1;dino_sprite[1][5][51] = 1;dino_sprite[1][5][52] = 1;dino_sprite[1][5][53] = 1;dino_sprite[1][5][54] = 1;dino_sprite[1][5][55] = 1;dino_sprite[1][5][56] = 1;dino_sprite[1][5][57] = 1;dino_sprite[1][5][58] = 1;dino_sprite[1][5][59] = 1;dino_sprite[1][5][60] = 1;dino_sprite[1][5][61] = 1;dino_sprite[1][5][62] = 1;dino_sprite[1][6][35] = 1;dino_sprite[1][6][36] = 1;dino_sprite[1][6][37] = 1;dino_sprite[1][6][38] = 1;dino_sprite[1][6][39] = 1;dino_sprite[1][6][40] = 1;dino_sprite[1][6][41] = 1;dino_sprite[1][6][42] = 1;dino_sprite[1][6][43] = 1;dino_sprite[1][6][44] = 1;dino_sprite[1][6][45] = 1;dino_sprite[1][6][46] = 1;dino_sprite[1][6][47] = 1;dino_sprite[1][6][48] = 1;dino_sprite[1][6][49] = 1;dino_sprite[1][6][50] = 1;dino_sprite[1][6][51] = 1;dino_sprite[1][6][52] = 1;dino_sprite[1][6][53] = 1;dino_sprite[1][6][54] = 1;dino_sprite[1][6][55] = 1;dino_sprite[1][6][56] = 1;dino_sprite[1][6][57] = 1;dino_sprite[1][6][58] = 1;dino_sprite[1][6][59] = 1;dino_sprite[1][6][60] = 1;dino_sprite[1][6][61] = 1;dino_sprite[1][6][62] = 1;dino_sprite[1][7][35] = 1;dino_sprite[1][7][36] = 1;dino_sprite[1][7][37] = 1;dino_sprite[1][7][38] = 1;dino_sprite[1][7][39] = 1;dino_sprite[1][7][40] = 1;dino_sprite[1][7][41] = 1;dino_sprite[1][7][42] = 1;dino_sprite[1][7][43] = 1;dino_sprite[1][7][44] = 1;dino_sprite[1][7][45] = 1;dino_sprite[1][7][46] = 1;dino_sprite[1][7][47] = 1;dino_sprite[1][7][48] = 1;dino_sprite[1][7][49] = 1;dino_sprite[1][7][50] = 1;dino_sprite[1][7][51] = 1;dino_sprite[1][7][52] = 1;dino_sprite[1][7][53] = 1;dino_sprite[1][7][54] = 1;dino_sprite[1][7][55] = 1;dino_sprite[1][7][56] = 1;dino_sprite[1][7][57] = 1;dino_sprite[1][7][58] = 1;dino_sprite[1][7][59] = 1;dino_sprite[1][7][60] = 1;dino_sprite[1][7][61] = 1;dino_sprite[1][7][62] = 1;dino_sprite[1][7][63] = 1;dino_sprite[1][7][64] = 1;dino_sprite[1][7][65] = 1;dino_sprite[1][7][66] = 1;dino_sprite[1][7][67] = 1;dino_sprite[1][8][44] = 1;dino_sprite[1][8][45] = 1;dino_sprite[1][8][46] = 1;dino_sprite[1][8][47] = 1;dino_sprite[1][8][48] = 1;dino_sprite[1][8][49] = 1;dino_sprite[1][8][50] = 1;dino_sprite[1][8][51] = 1;dino_sprite[1][8][52] = 1;dino_sprite[1][8][53] = 1;dino_sprite[1][8][54] = 1;dino_sprite[1][8][55] = 1;dino_sprite[1][8][56] = 1;dino_sprite[1][8][57] = 1;dino_sprite[1][8][58] = 1;dino_sprite[1][8][59] = 1;dino_sprite[1][8][60] = 1;dino_sprite[1][8][61] = 1;dino_sprite[1][8][62] = 1;dino_sprite[1][8][63] = 1;dino_sprite[1][8][64] = 1;dino_sprite[1][8][65] = 1;dino_sprite[1][8][66] = 1;dino_sprite[1][8][67] = 1;dino_sprite[1][9][44] = 1;dino_sprite[1][9][45] = 1;dino_sprite[1][9][46] = 1;dino_sprite[1][9][47] = 1;dino_sprite[1][9][48] = 1;dino_sprite[1][9][49] = 1;dino_sprite[1][9][50] = 1;dino_sprite[1][9][51] = 1;dino_sprite[1][9][52] = 1;dino_sprite[1][9][53] = 1;dino_sprite[1][9][54] = 1;dino_sprite[1][9][55] = 1;dino_sprite[1][9][56] = 1;dino_sprite[1][9][57] = 1;dino_sprite[1][9][58] = 1;dino_sprite[1][9][59] = 1;dino_sprite[1][9][60] = 1;dino_sprite[1][9][61] = 1;dino_sprite[1][9][62] = 1;dino_sprite[1][9][63] = 1;dino_sprite[1][9][64] = 1;dino_sprite[1][9][65] = 1;dino_sprite[1][9][66] = 1;dino_sprite[1][9][67] = 1;dino_sprite[1][10][44] = 1;dino_sprite[1][10][45] = 1;dino_sprite[1][10][46] = 1;dino_sprite[1][10][47] = 1;dino_sprite[1][10][48] = 1;dino_sprite[1][10][49] = 1;dino_sprite[1][10][50] = 1;dino_sprite[1][10][51] = 1;dino_sprite[1][10][52] = 1;dino_sprite[1][10][53] = 1;dino_sprite[1][10][54] = 1;dino_sprite[1][10][55] = 1;dino_sprite[1][10][56] = 1;dino_sprite[1][10][57] = 1;dino_sprite[1][10][58] = 1;dino_sprite[1][10][59] = 1;dino_sprite[1][10][60] = 1;dino_sprite[1][10][61] = 1;dino_sprite[1][10][62] = 1;dino_sprite[1][10][63] = 1;dino_sprite[1][10][64] = 1;dino_sprite[1][10][65] = 1;dino_sprite[1][10][66] = 1;dino_sprite[1][10][67] = 1;dino_sprite[1][11][44] = 1;dino_sprite[1][11][45] = 1;dino_sprite[1][11][46] = 1;dino_sprite[1][11][47] = 1;dino_sprite[1][11][48] = 1;dino_sprite[1][11][49] = 1;dino_sprite[1][11][50] = 1;dino_sprite[1][11][51] = 1;dino_sprite[1][11][52] = 1;dino_sprite[1][11][53] = 1;dino_sprite[1][11][54] = 1;dino_sprite[1][11][55] = 1;dino_sprite[1][11][56] = 1;dino_sprite[1][11][57] = 1;dino_sprite[1][11][58] = 1;dino_sprite[1][11][59] = 1;dino_sprite[1][11][60] = 1;dino_sprite[1][11][61] = 1;dino_sprite[1][11][62] = 1;dino_sprite[1][11][63] = 1;dino_sprite[1][11][64] = 1;dino_sprite[1][11][65] = 1;dino_sprite[1][11][66] = 1;dino_sprite[1][11][67] = 1;dino_sprite[1][12][49] = 1;dino_sprite[1][12][50] = 1;dino_sprite[1][12][51] = 1;dino_sprite[1][12][52] = 1;dino_sprite[1][12][53] = 1;dino_sprite[1][12][54] = 1;dino_sprite[1][12][55] = 1;dino_sprite[1][12][56] = 1;dino_sprite[1][12][57] = 1;dino_sprite[1][12][58] = 1;dino_sprite[1][12][59] = 1;dino_sprite[1][12][60] = 1;dino_sprite[1][12][61] = 1;dino_sprite[1][12][62] = 1;dino_sprite[1][12][63] = 1;dino_sprite[1][12][64] = 1;dino_sprite[1][12][65] = 1;dino_sprite[1][12][66] = 1;dino_sprite[1][12][67] = 1;dino_sprite[1][12][68] = 1;dino_sprite[1][12][69] = 1;dino_sprite[1][12][70] = 1;dino_sprite[1][12][71] = 1;dino_sprite[1][12][72] = 1;dino_sprite[1][13][49] = 1;dino_sprite[1][13][50] = 1;dino_sprite[1][13][51] = 1;dino_sprite[1][13][52] = 1;dino_sprite[1][13][53] = 1;dino_sprite[1][13][54] = 1;dino_sprite[1][13][55] = 1;dino_sprite[1][13][56] = 1;dino_sprite[1][13][57] = 1;dino_sprite[1][13][58] = 1;dino_sprite[1][13][59] = 1;dino_sprite[1][13][60] = 1;dino_sprite[1][13][61] = 1;dino_sprite[1][13][62] = 1;dino_sprite[1][13][63] = 1;dino_sprite[1][13][64] = 1;dino_sprite[1][13][65] = 1;dino_sprite[1][13][66] = 1;dino_sprite[1][13][67] = 1;dino_sprite[1][13][68] = 1;dino_sprite[1][13][69] = 1;dino_sprite[1][13][70] = 1;dino_sprite[1][13][71] = 1;dino_sprite[1][13][72] = 1;dino_sprite[1][14][49] = 1;dino_sprite[1][14][50] = 1;dino_sprite[1][14][51] = 1;dino_sprite[1][14][52] = 1;dino_sprite[1][14][53] = 1;dino_sprite[1][14][54] = 1;dino_sprite[1][14][55] = 1;dino_sprite[1][14][56] = 1;dino_sprite[1][14][57] = 1;dino_sprite[1][14][58] = 1;dino_sprite[1][14][59] = 1;dino_sprite[1][14][60] = 1;dino_sprite[1][14][61] = 1;dino_sprite[1][14][62] = 1;dino_sprite[1][14][63] = 1;dino_sprite[1][14][64] = 1;dino_sprite[1][14][65] = 1;dino_sprite[1][14][66] = 1;dino_sprite[1][14][67] = 1;dino_sprite[1][14][68] = 1;dino_sprite[1][14][69] = 1;dino_sprite[1][14][70] = 1;dino_sprite[1][14][71] = 1;dino_sprite[1][14][72] = 1;dino_sprite[1][15][49] = 1;dino_sprite[1][15][50] = 1;dino_sprite[1][15][51] = 1;dino_sprite[1][15][52] = 1;dino_sprite[1][15][53] = 1;dino_sprite[1][15][54] = 1;dino_sprite[1][15][55] = 1;dino_sprite[1][15][56] = 1;dino_sprite[1][15][57] = 1;dino_sprite[1][15][58] = 1;dino_sprite[1][15][59] = 1;dino_sprite[1][15][60] = 1;dino_sprite[1][15][61] = 1;dino_sprite[1][15][62] = 1;dino_sprite[1][15][63] = 1;dino_sprite[1][15][64] = 1;dino_sprite[1][15][65] = 1;dino_sprite[1][15][66] = 1;dino_sprite[1][15][67] = 1;dino_sprite[1][15][68] = 1;dino_sprite[1][15][69] = 1;dino_sprite[1][15][70] = 1;dino_sprite[1][15][71] = 1;dino_sprite[1][15][72] = 1;dino_sprite[1][16][49] = 1;dino_sprite[1][16][50] = 1;dino_sprite[1][16][51] = 1;dino_sprite[1][16][52] = 1;dino_sprite[1][16][53] = 1;dino_sprite[1][16][54] = 1;dino_sprite[1][16][55] = 1;dino_sprite[1][16][56] = 1;dino_sprite[1][16][57] = 1;dino_sprite[1][16][58] = 1;dino_sprite[1][16][59] = 1;dino_sprite[1][16][60] = 1;dino_sprite[1][16][61] = 1;dino_sprite[1][16][62] = 1;dino_sprite[1][16][63] = 1;dino_sprite[1][16][64] = 1;dino_sprite[1][16][65] = 1;dino_sprite[1][16][66] = 1;dino_sprite[1][16][67] = 1;dino_sprite[1][16][68] = 1;dino_sprite[1][16][69] = 1;dino_sprite[1][16][70] = 1;dino_sprite[1][16][71] = 1;dino_sprite[1][16][72] = 1;dino_sprite[1][17][54] = 1;dino_sprite[1][17][55] = 1;dino_sprite[1][17][56] = 1;dino_sprite[1][17][57] = 1;dino_sprite[1][17][58] = 1;dino_sprite[1][17][59] = 1;dino_sprite[1][17][60] = 1;dino_sprite[1][17][61] = 1;dino_sprite[1][17][62] = 1;dino_sprite[1][17][63] = 1;dino_sprite[1][17][64] = 1;dino_sprite[1][17][65] = 1;dino_sprite[1][17][66] = 1;dino_sprite[1][17][67] = 1;dino_sprite[1][17][68] = 1;dino_sprite[1][17][69] = 1;dino_sprite[1][17][70] = 1;dino_sprite[1][17][71] = 1;dino_sprite[1][17][72] = 1;dino_sprite[1][17][73] = 1;dino_sprite[1][17][74] = 1;dino_sprite[1][17][75] = 1;dino_sprite[1][17][76] = 1;dino_sprite[1][17][77] = 1;dino_sprite[1][18][54] = 1;dino_sprite[1][18][55] = 1;dino_sprite[1][18][56] = 1;dino_sprite[1][18][57] = 1;dino_sprite[1][18][58] = 1;dino_sprite[1][18][59] = 1;dino_sprite[1][18][60] = 1;dino_sprite[1][18][61] = 1;dino_sprite[1][18][62] = 1;dino_sprite[1][18][63] = 1;dino_sprite[1][18][64] = 1;dino_sprite[1][18][65] = 1;dino_sprite[1][18][66] = 1;dino_sprite[1][18][67] = 1;dino_sprite[1][18][68] = 1;dino_sprite[1][18][69] = 1;dino_sprite[1][18][70] = 1;dino_sprite[1][18][71] = 1;dino_sprite[1][18][72] = 1;dino_sprite[1][18][73] = 1;dino_sprite[1][18][74] = 1;dino_sprite[1][18][75] = 1;dino_sprite[1][18][76] = 1;dino_sprite[1][18][77] = 1;dino_sprite[1][19][54] = 1;dino_sprite[1][19][55] = 1;dino_sprite[1][19][56] = 1;dino_sprite[1][19][57] = 1;dino_sprite[1][19][58] = 1;dino_sprite[1][19][59] = 1;dino_sprite[1][19][60] = 1;dino_sprite[1][19][61] = 1;dino_sprite[1][19][62] = 1;dino_sprite[1][19][63] = 1;dino_sprite[1][19][64] = 1;dino_sprite[1][19][65] = 1;dino_sprite[1][19][66] = 1;dino_sprite[1][19][67] = 1;dino_sprite[1][19][68] = 1;dino_sprite[1][19][69] = 1;dino_sprite[1][19][70] = 1;dino_sprite[1][19][71] = 1;dino_sprite[1][19][72] = 1;dino_sprite[1][19][73] = 1;dino_sprite[1][19][74] = 1;dino_sprite[1][19][75] = 1;dino_sprite[1][19][76] = 1;dino_sprite[1][19][77] = 1;dino_sprite[1][20][54] = 1;dino_sprite[1][20][55] = 1;dino_sprite[1][20][56] = 1;dino_sprite[1][20][57] = 1;dino_sprite[1][20][58] = 1;dino_sprite[1][20][59] = 1;dino_sprite[1][20][60] = 1;dino_sprite[1][20][61] = 1;dino_sprite[1][20][62] = 1;dino_sprite[1][20][63] = 1;dino_sprite[1][20][64] = 1;dino_sprite[1][20][65] = 1;dino_sprite[1][20][66] = 1;dino_sprite[1][20][67] = 1;dino_sprite[1][20][68] = 1;dino_sprite[1][20][69] = 1;dino_sprite[1][20][70] = 1;dino_sprite[1][20][71] = 1;dino_sprite[1][20][72] = 1;dino_sprite[1][20][73] = 1;dino_sprite[1][20][74] = 1;dino_sprite[1][20][75] = 1;dino_sprite[1][20][76] = 1;dino_sprite[1][20][77] = 1;dino_sprite[1][21][54] = 1;dino_sprite[1][21][55] = 1;dino_sprite[1][21][56] = 1;dino_sprite[1][21][57] = 1;dino_sprite[1][21][58] = 1;dino_sprite[1][21][59] = 1;dino_sprite[1][21][60] = 1;dino_sprite[1][21][61] = 1;dino_sprite[1][21][62] = 1;dino_sprite[1][21][63] = 1;dino_sprite[1][21][64] = 1;dino_sprite[1][21][65] = 1;dino_sprite[1][21][66] = 1;dino_sprite[1][21][67] = 1;dino_sprite[1][21][68] = 1;dino_sprite[1][21][69] = 1;dino_sprite[1][21][70] = 1;dino_sprite[1][21][71] = 1;dino_sprite[1][21][72] = 1;dino_sprite[1][21][73] = 1;dino_sprite[1][21][74] = 1;dino_sprite[1][21][75] = 1;dino_sprite[1][21][76] = 1;dino_sprite[1][21][77] = 1;dino_sprite[1][22][54] = 1;dino_sprite[1][22][55] = 1;dino_sprite[1][22][56] = 1;dino_sprite[1][22][57] = 1;dino_sprite[1][22][58] = 1;dino_sprite[1][22][59] = 1;dino_sprite[1][22][60] = 1;dino_sprite[1][22][61] = 1;dino_sprite[1][22][62] = 1;dino_sprite[1][22][63] = 1;dino_sprite[1][22][64] = 1;dino_sprite[1][22][65] = 1;dino_sprite[1][22][66] = 1;dino_sprite[1][22][67] = 1;dino_sprite[1][22][68] = 1;dino_sprite[1][22][69] = 1;dino_sprite[1][22][70] = 1;dino_sprite[1][22][71] = 1;dino_sprite[1][22][72] = 1;dino_sprite[1][22][73] = 1;dino_sprite[1][22][74] = 1;dino_sprite[1][22][75] = 1;dino_sprite[1][22][76] = 1;dino_sprite[1][22][77] = 1;dino_sprite[1][22][78] = 1;dino_sprite[1][22][79] = 1;dino_sprite[1][22][80] = 1;dino_sprite[1][22][81] = 1;dino_sprite[1][23][54] = 1;dino_sprite[1][23][55] = 1;dino_sprite[1][23][56] = 1;dino_sprite[1][23][57] = 1;dino_sprite[1][23][58] = 1;dino_sprite[1][23][59] = 1;dino_sprite[1][23][60] = 1;dino_sprite[1][23][61] = 1;dino_sprite[1][23][62] = 1;dino_sprite[1][23][63] = 1;dino_sprite[1][23][64] = 1;dino_sprite[1][23][65] = 1;dino_sprite[1][23][66] = 1;dino_sprite[1][23][67] = 1;dino_sprite[1][23][68] = 1;dino_sprite[1][23][69] = 1;dino_sprite[1][23][70] = 1;dino_sprite[1][23][71] = 1;dino_sprite[1][23][72] = 1;dino_sprite[1][23][73] = 1;dino_sprite[1][23][74] = 1;dino_sprite[1][23][75] = 1;dino_sprite[1][23][76] = 1;dino_sprite[1][23][77] = 1;dino_sprite[1][23][78] = 1;dino_sprite[1][23][79] = 1;dino_sprite[1][23][80] = 1;dino_sprite[1][23][81] = 1;dino_sprite[1][24][54] = 1;dino_sprite[1][24][55] = 1;dino_sprite[1][24][56] = 1;dino_sprite[1][24][57] = 1;dino_sprite[1][24][58] = 1;dino_sprite[1][24][59] = 1;dino_sprite[1][24][60] = 1;dino_sprite[1][24][61] = 1;dino_sprite[1][24][62] = 1;dino_sprite[1][24][63] = 1;dino_sprite[1][24][64] = 1;dino_sprite[1][24][65] = 1;dino_sprite[1][24][66] = 1;dino_sprite[1][24][67] = 1;dino_sprite[1][24][68] = 1;dino_sprite[1][24][69] = 1;dino_sprite[1][24][70] = 1;dino_sprite[1][24][71] = 1;dino_sprite[1][24][72] = 1;dino_sprite[1][24][73] = 1;dino_sprite[1][24][74] = 1;dino_sprite[1][24][75] = 1;dino_sprite[1][24][76] = 1;dino_sprite[1][24][77] = 1;dino_sprite[1][24][78] = 1;dino_sprite[1][24][79] = 1;dino_sprite[1][24][80] = 1;dino_sprite[1][24][81] = 1;dino_sprite[1][25][54] = 1;dino_sprite[1][25][55] = 1;dino_sprite[1][25][56] = 1;dino_sprite[1][25][57] = 1;dino_sprite[1][25][58] = 1;dino_sprite[1][25][59] = 1;dino_sprite[1][25][60] = 1;dino_sprite[1][25][61] = 1;dino_sprite[1][25][62] = 1;dino_sprite[1][25][63] = 1;dino_sprite[1][25][64] = 1;dino_sprite[1][25][65] = 1;dino_sprite[1][25][66] = 1;dino_sprite[1][25][67] = 1;dino_sprite[1][25][68] = 1;dino_sprite[1][25][69] = 1;dino_sprite[1][25][70] = 1;dino_sprite[1][25][71] = 1;dino_sprite[1][25][72] = 1;dino_sprite[1][25][73] = 1;dino_sprite[1][25][74] = 1;dino_sprite[1][25][75] = 1;dino_sprite[1][25][76] = 1;dino_sprite[1][25][77] = 1;dino_sprite[1][25][78] = 1;dino_sprite[1][25][79] = 1;dino_sprite[1][25][80] = 1;dino_sprite[1][25][81] = 1;dino_sprite[1][26][49] = 1;dino_sprite[1][26][50] = 1;dino_sprite[1][26][51] = 1;dino_sprite[1][26][52] = 1;dino_sprite[1][26][53] = 1;dino_sprite[1][26][54] = 1;dino_sprite[1][26][55] = 1;dino_sprite[1][26][56] = 1;dino_sprite[1][26][57] = 1;dino_sprite[1][26][58] = 1;dino_sprite[1][26][59] = 1;dino_sprite[1][26][60] = 1;dino_sprite[1][26][61] = 1;dino_sprite[1][26][62] = 1;dino_sprite[1][26][63] = 1;dino_sprite[1][26][64] = 1;dino_sprite[1][26][65] = 1;dino_sprite[1][26][66] = 1;dino_sprite[1][26][67] = 1;dino_sprite[1][26][68] = 1;dino_sprite[1][26][69] = 1;dino_sprite[1][26][70] = 1;dino_sprite[1][26][71] = 1;dino_sprite[1][26][72] = 1;dino_sprite[1][26][73] = 1;dino_sprite[1][26][74] = 1;dino_sprite[1][26][75] = 1;dino_sprite[1][26][76] = 1;dino_sprite[1][26][77] = 1;dino_sprite[1][26][78] = 1;dino_sprite[1][26][79] = 1;dino_sprite[1][26][80] = 1;dino_sprite[1][26][81] = 1;dino_sprite[1][26][82] = 1;dino_sprite[1][26][83] = 1;dino_sprite[1][26][84] = 1;dino_sprite[1][26][85] = 1;dino_sprite[1][26][86] = 1;dino_sprite[1][26][87] = 1;dino_sprite[1][26][88] = 1;dino_sprite[1][26][89] = 1;dino_sprite[1][26][90] = 1;dino_sprite[1][26][91] = 1;dino_sprite[1][26][92] = 1;dino_sprite[1][27][49] = 1;dino_sprite[1][27][50] = 1;dino_sprite[1][27][51] = 1;dino_sprite[1][27][52] = 1;dino_sprite[1][27][53] = 1;dino_sprite[1][27][54] = 1;dino_sprite[1][27][55] = 1;dino_sprite[1][27][56] = 1;dino_sprite[1][27][57] = 1;dino_sprite[1][27][58] = 1;dino_sprite[1][27][59] = 1;dino_sprite[1][27][60] = 1;dino_sprite[1][27][61] = 1;dino_sprite[1][27][62] = 1;dino_sprite[1][27][63] = 1;dino_sprite[1][27][64] = 1;dino_sprite[1][27][65] = 1;dino_sprite[1][27][66] = 1;dino_sprite[1][27][67] = 1;dino_sprite[1][27][68] = 1;dino_sprite[1][27][69] = 1;dino_sprite[1][27][70] = 1;dino_sprite[1][27][71] = 1;dino_sprite[1][27][72] = 1;dino_sprite[1][27][73] = 1;dino_sprite[1][27][74] = 1;dino_sprite[1][27][75] = 1;dino_sprite[1][27][76] = 1;dino_sprite[1][27][77] = 1;dino_sprite[1][27][78] = 1;dino_sprite[1][27][79] = 1;dino_sprite[1][27][80] = 1;dino_sprite[1][27][81] = 1;dino_sprite[1][27][82] = 1;dino_sprite[1][27][83] = 1;dino_sprite[1][27][84] = 1;dino_sprite[1][27][85] = 1;dino_sprite[1][27][86] = 1;dino_sprite[1][27][87] = 1;dino_sprite[1][27][88] = 1;dino_sprite[1][27][89] = 1;dino_sprite[1][27][90] = 1;dino_sprite[1][27][91] = 1;dino_sprite[1][27][92] = 1;dino_sprite[1][28][49] = 1;dino_sprite[1][28][50] = 1;dino_sprite[1][28][51] = 1;dino_sprite[1][28][52] = 1;dino_sprite[1][28][53] = 1;dino_sprite[1][28][54] = 1;dino_sprite[1][28][55] = 1;dino_sprite[1][28][56] = 1;dino_sprite[1][28][57] = 1;dino_sprite[1][28][58] = 1;dino_sprite[1][28][59] = 1;dino_sprite[1][28][60] = 1;dino_sprite[1][28][61] = 1;dino_sprite[1][28][62] = 1;dino_sprite[1][28][63] = 1;dino_sprite[1][28][64] = 1;dino_sprite[1][28][65] = 1;dino_sprite[1][28][66] = 1;dino_sprite[1][28][67] = 1;dino_sprite[1][28][68] = 1;dino_sprite[1][28][69] = 1;dino_sprite[1][28][70] = 1;dino_sprite[1][28][71] = 1;dino_sprite[1][28][72] = 1;dino_sprite[1][28][73] = 1;dino_sprite[1][28][74] = 1;dino_sprite[1][28][75] = 1;dino_sprite[1][28][76] = 1;dino_sprite[1][28][77] = 1;dino_sprite[1][28][78] = 1;dino_sprite[1][28][79] = 1;dino_sprite[1][28][80] = 1;dino_sprite[1][28][81] = 1;dino_sprite[1][28][82] = 1;dino_sprite[1][28][83] = 1;dino_sprite[1][28][84] = 1;dino_sprite[1][28][85] = 1;dino_sprite[1][28][86] = 1;dino_sprite[1][28][87] = 1;dino_sprite[1][28][88] = 1;dino_sprite[1][28][89] = 1;dino_sprite[1][28][90] = 1;dino_sprite[1][28][91] = 1;dino_sprite[1][28][92] = 1;dino_sprite[1][29][49] = 1;dino_sprite[1][29][50] = 1;dino_sprite[1][29][51] = 1;dino_sprite[1][29][52] = 1;dino_sprite[1][29][53] = 1;dino_sprite[1][29][54] = 1;dino_sprite[1][29][55] = 1;dino_sprite[1][29][56] = 1;dino_sprite[1][29][57] = 1;dino_sprite[1][29][58] = 1;dino_sprite[1][29][59] = 1;dino_sprite[1][29][60] = 1;dino_sprite[1][29][61] = 1;dino_sprite[1][29][62] = 1;dino_sprite[1][29][63] = 1;dino_sprite[1][29][64] = 1;dino_sprite[1][29][65] = 1;dino_sprite[1][29][66] = 1;dino_sprite[1][29][67] = 1;dino_sprite[1][29][68] = 1;dino_sprite[1][29][69] = 1;dino_sprite[1][29][70] = 1;dino_sprite[1][29][71] = 1;dino_sprite[1][29][72] = 1;dino_sprite[1][29][73] = 1;dino_sprite[1][29][74] = 1;dino_sprite[1][29][75] = 1;dino_sprite[1][29][76] = 1;dino_sprite[1][29][77] = 1;dino_sprite[1][29][78] = 1;dino_sprite[1][29][79] = 1;dino_sprite[1][29][80] = 1;dino_sprite[1][29][81] = 1;dino_sprite[1][29][82] = 1;dino_sprite[1][29][83] = 1;dino_sprite[1][29][84] = 1;dino_sprite[1][29][85] = 1;dino_sprite[1][29][86] = 1;dino_sprite[1][29][87] = 1;dino_sprite[1][29][88] = 1;dino_sprite[1][29][89] = 1;dino_sprite[1][29][90] = 1;dino_sprite[1][29][91] = 1;dino_sprite[1][29][92] = 1;dino_sprite[1][30][49] = 1;dino_sprite[1][30][50] = 1;dino_sprite[1][30][51] = 1;dino_sprite[1][30][52] = 1;dino_sprite[1][30][53] = 1;dino_sprite[1][30][54] = 1;dino_sprite[1][30][55] = 1;dino_sprite[1][30][56] = 1;dino_sprite[1][30][57] = 1;dino_sprite[1][30][58] = 1;dino_sprite[1][30][59] = 1;dino_sprite[1][30][60] = 1;dino_sprite[1][30][61] = 1;dino_sprite[1][30][62] = 1;dino_sprite[1][30][63] = 1;dino_sprite[1][30][64] = 1;dino_sprite[1][30][65] = 1;dino_sprite[1][30][66] = 1;dino_sprite[1][30][67] = 1;dino_sprite[1][30][68] = 1;dino_sprite[1][30][69] = 1;dino_sprite[1][30][70] = 1;dino_sprite[1][30][71] = 1;dino_sprite[1][30][72] = 1;dino_sprite[1][30][73] = 1;dino_sprite[1][30][74] = 1;dino_sprite[1][30][75] = 1;dino_sprite[1][30][76] = 1;dino_sprite[1][30][77] = 1;dino_sprite[1][30][78] = 1;dino_sprite[1][30][79] = 1;dino_sprite[1][30][80] = 1;dino_sprite[1][30][81] = 1;dino_sprite[1][30][82] = 1;dino_sprite[1][30][83] = 1;dino_sprite[1][30][84] = 1;dino_sprite[1][30][85] = 1;dino_sprite[1][30][86] = 1;dino_sprite[1][30][87] = 1;dino_sprite[1][30][88] = 1;dino_sprite[1][30][89] = 1;dino_sprite[1][30][90] = 1;dino_sprite[1][30][91] = 1;dino_sprite[1][30][92] = 1;dino_sprite[1][31][44] = 1;dino_sprite[1][31][45] = 1;dino_sprite[1][31][46] = 1;dino_sprite[1][31][47] = 1;dino_sprite[1][31][48] = 1;dino_sprite[1][31][49] = 1;dino_sprite[1][31][50] = 1;dino_sprite[1][31][51] = 1;dino_sprite[1][31][52] = 1;dino_sprite[1][31][53] = 1;dino_sprite[1][31][54] = 1;dino_sprite[1][31][55] = 1;dino_sprite[1][31][56] = 1;dino_sprite[1][31][57] = 1;dino_sprite[1][31][58] = 1;dino_sprite[1][31][59] = 1;dino_sprite[1][31][60] = 1;dino_sprite[1][31][61] = 1;dino_sprite[1][31][62] = 1;dino_sprite[1][31][63] = 1;dino_sprite[1][31][64] = 1;dino_sprite[1][31][65] = 1;dino_sprite[1][31][66] = 1;dino_sprite[1][31][67] = 1;dino_sprite[1][31][68] = 1;dino_sprite[1][31][69] = 1;dino_sprite[1][31][70] = 1;dino_sprite[1][31][71] = 1;dino_sprite[1][31][72] = 1;dino_sprite[1][31][73] = 1;dino_sprite[1][31][74] = 1;dino_sprite[1][31][75] = 1;dino_sprite[1][31][76] = 1;dino_sprite[1][31][77] = 1;dino_sprite[1][31][78] = 1;dino_sprite[1][31][79] = 1;dino_sprite[1][31][80] = 1;dino_sprite[1][31][81] = 1;dino_sprite[1][31][82] = 1;dino_sprite[1][31][83] = 1;dino_sprite[1][31][84] = 1;dino_sprite[1][31][85] = 1;dino_sprite[1][31][86] = 1;dino_sprite[1][31][87] = 1;dino_sprite[1][31][88] = 1;dino_sprite[1][31][89] = 1;dino_sprite[1][31][90] = 1;dino_sprite[1][31][91] = 1;dino_sprite[1][31][92] = 1;dino_sprite[1][32][44] = 1;dino_sprite[1][32][45] = 1;dino_sprite[1][32][46] = 1;dino_sprite[1][32][47] = 1;dino_sprite[1][32][48] = 1;dino_sprite[1][32][49] = 1;dino_sprite[1][32][50] = 1;dino_sprite[1][32][51] = 1;dino_sprite[1][32][52] = 1;dino_sprite[1][32][53] = 1;dino_sprite[1][32][54] = 1;dino_sprite[1][32][55] = 1;dino_sprite[1][32][56] = 1;dino_sprite[1][32][57] = 1;dino_sprite[1][32][58] = 1;dino_sprite[1][32][59] = 1;dino_sprite[1][32][60] = 1;dino_sprite[1][32][61] = 1;dino_sprite[1][32][62] = 1;dino_sprite[1][32][63] = 1;dino_sprite[1][32][64] = 1;dino_sprite[1][32][65] = 1;dino_sprite[1][32][66] = 1;dino_sprite[1][32][67] = 1;dino_sprite[1][32][68] = 1;dino_sprite[1][32][69] = 1;dino_sprite[1][32][70] = 1;dino_sprite[1][32][71] = 1;dino_sprite[1][32][72] = 1;dino_sprite[1][32][73] = 1;dino_sprite[1][32][74] = 1;dino_sprite[1][32][75] = 1;dino_sprite[1][32][76] = 1;dino_sprite[1][32][77] = 1;dino_sprite[1][32][78] = 1;dino_sprite[1][32][79] = 1;dino_sprite[1][32][80] = 1;dino_sprite[1][32][81] = 1;dino_sprite[1][32][82] = 1;dino_sprite[1][32][83] = 1;dino_sprite[1][32][84] = 1;dino_sprite[1][32][85] = 1;dino_sprite[1][32][86] = 1;dino_sprite[1][32][88] = 1;dino_sprite[1][32][89] = 1;dino_sprite[1][32][90] = 1;dino_sprite[1][32][91] = 1;dino_sprite[1][32][92] = 1;dino_sprite[1][33][44] = 1;dino_sprite[1][33][45] = 1;dino_sprite[1][33][46] = 1;dino_sprite[1][33][47] = 1;dino_sprite[1][33][48] = 1;dino_sprite[1][33][49] = 1;dino_sprite[1][33][50] = 1;dino_sprite[1][33][51] = 1;dino_sprite[1][33][52] = 1;dino_sprite[1][33][53] = 1;dino_sprite[1][33][54] = 1;dino_sprite[1][33][55] = 1;dino_sprite[1][33][56] = 1;dino_sprite[1][33][57] = 1;dino_sprite[1][33][58] = 1;dino_sprite[1][33][59] = 1;dino_sprite[1][33][60] = 1;dino_sprite[1][33][61] = 1;dino_sprite[1][33][62] = 1;dino_sprite[1][33][63] = 1;dino_sprite[1][33][64] = 1;dino_sprite[1][33][65] = 1;dino_sprite[1][33][66] = 1;dino_sprite[1][33][67] = 1;dino_sprite[1][33][68] = 1;dino_sprite[1][33][69] = 1;dino_sprite[1][33][70] = 1;dino_sprite[1][33][71] = 1;dino_sprite[1][33][72] = 1;dino_sprite[1][33][73] = 1;dino_sprite[1][33][74] = 1;dino_sprite[1][33][75] = 1;dino_sprite[1][33][76] = 1;dino_sprite[1][33][77] = 1;dino_sprite[1][33][78] = 1;dino_sprite[1][33][79] = 1;dino_sprite[1][33][80] = 1;dino_sprite[1][33][81] = 1;dino_sprite[1][33][82] = 1;dino_sprite[1][33][83] = 1;dino_sprite[1][33][84] = 1;dino_sprite[1][33][85] = 1;dino_sprite[1][33][86] = 1;dino_sprite[1][33][88] = 1;dino_sprite[1][33][89] = 1;dino_sprite[1][33][90] = 1;dino_sprite[1][33][91] = 1;dino_sprite[1][33][92] = 1;dino_sprite[1][34][44] = 1;dino_sprite[1][34][45] = 1;dino_sprite[1][34][46] = 1;dino_sprite[1][34][47] = 1;dino_sprite[1][34][48] = 1;dino_sprite[1][34][49] = 1;dino_sprite[1][34][50] = 1;dino_sprite[1][34][51] = 1;dino_sprite[1][34][52] = 1;dino_sprite[1][34][53] = 1;dino_sprite[1][34][54] = 1;dino_sprite[1][34][55] = 1;dino_sprite[1][34][56] = 1;dino_sprite[1][34][57] = 1;dino_sprite[1][34][58] = 1;dino_sprite[1][34][59] = 1;dino_sprite[1][34][60] = 1;dino_sprite[1][34][61] = 1;dino_sprite[1][34][62] = 1;dino_sprite[1][34][63] = 1;dino_sprite[1][34][64] = 1;dino_sprite[1][34][65] = 1;dino_sprite[1][34][66] = 1;dino_sprite[1][34][67] = 1;dino_sprite[1][34][68] = 1;dino_sprite[1][34][69] = 1;dino_sprite[1][34][70] = 1;dino_sprite[1][34][71] = 1;dino_sprite[1][34][72] = 1;dino_sprite[1][34][73] = 1;dino_sprite[1][34][74] = 1;dino_sprite[1][34][75] = 1;dino_sprite[1][34][76] = 1;dino_sprite[1][34][77] = 1;dino_sprite[1][34][78] = 1;dino_sprite[1][34][79] = 1;dino_sprite[1][34][80] = 1;dino_sprite[1][34][81] = 1;dino_sprite[1][34][82] = 1;dino_sprite[1][34][83] = 1;dino_sprite[1][34][84] = 1;dino_sprite[1][34][85] = 1;dino_sprite[1][34][86] = 1;dino_sprite[1][34][88] = 1;dino_sprite[1][34][89] = 1;dino_sprite[1][34][90] = 1;dino_sprite[1][34][91] = 1;dino_sprite[1][34][92] = 1;dino_sprite[1][35][44] = 1;dino_sprite[1][35][45] = 1;dino_sprite[1][35][46] = 1;dino_sprite[1][35][47] = 1;dino_sprite[1][35][48] = 1;dino_sprite[1][35][49] = 1;dino_sprite[1][35][50] = 1;dino_sprite[1][35][51] = 1;dino_sprite[1][35][52] = 1;dino_sprite[1][35][53] = 1;dino_sprite[1][35][54] = 1;dino_sprite[1][35][55] = 1;dino_sprite[1][35][56] = 1;dino_sprite[1][35][57] = 1;dino_sprite[1][35][58] = 1;dino_sprite[1][35][59] = 1;dino_sprite[1][35][60] = 1;dino_sprite[1][35][61] = 1;dino_sprite[1][35][62] = 1;dino_sprite[1][35][63] = 1;dino_sprite[1][35][64] = 1;dino_sprite[1][35][65] = 1;dino_sprite[1][35][66] = 1;dino_sprite[1][35][67] = 1;dino_sprite[1][35][68] = 1;dino_sprite[1][35][69] = 1;dino_sprite[1][35][70] = 1;dino_sprite[1][35][71] = 1;dino_sprite[1][35][72] = 1;dino_sprite[1][35][73] = 1;dino_sprite[1][35][74] = 1;dino_sprite[1][35][75] = 1;dino_sprite[1][35][76] = 1;dino_sprite[1][35][77] = 1;dino_sprite[1][35][78] = 1;dino_sprite[1][35][79] = 1;dino_sprite[1][35][80] = 1;dino_sprite[1][35][81] = 1;dino_sprite[1][35][82] = 1;dino_sprite[1][35][83] = 1;dino_sprite[1][35][84] = 1;dino_sprite[1][35][85] = 1;dino_sprite[1][35][86] = 1;dino_sprite[1][35][88] = 1;dino_sprite[1][35][89] = 1;dino_sprite[1][35][90] = 1;dino_sprite[1][35][91] = 1;dino_sprite[1][35][92] = 1;dino_sprite[1][36][44] = 1;dino_sprite[1][36][45] = 1;dino_sprite[1][36][46] = 1;dino_sprite[1][36][47] = 1;dino_sprite[1][36][48] = 1;dino_sprite[1][36][49] = 1;dino_sprite[1][36][50] = 1;dino_sprite[1][36][51] = 1;dino_sprite[1][36][52] = 1;dino_sprite[1][36][53] = 1;dino_sprite[1][36][54] = 1;dino_sprite[1][36][55] = 1;dino_sprite[1][36][56] = 1;dino_sprite[1][36][57] = 1;dino_sprite[1][36][58] = 1;dino_sprite[1][36][59] = 1;dino_sprite[1][36][60] = 1;dino_sprite[1][36][61] = 1;dino_sprite[1][36][62] = 1;dino_sprite[1][36][63] = 1;dino_sprite[1][36][64] = 1;dino_sprite[1][36][65] = 1;dino_sprite[1][36][66] = 1;dino_sprite[1][36][67] = 1;dino_sprite[1][36][68] = 1;dino_sprite[1][36][69] = 1;dino_sprite[1][36][70] = 1;dino_sprite[1][36][71] = 1;dino_sprite[1][36][72] = 1;dino_sprite[1][36][73] = 1;dino_sprite[1][36][74] = 1;dino_sprite[1][36][75] = 1;dino_sprite[1][36][76] = 1;dino_sprite[1][36][77] = 1;dino_sprite[1][36][78] = 1;dino_sprite[1][36][79] = 1;dino_sprite[1][36][80] = 1;dino_sprite[1][36][81] = 1;dino_sprite[1][36][82] = 1;dino_sprite[1][36][83] = 1;dino_sprite[1][36][84] = 1;dino_sprite[1][36][85] = 1;dino_sprite[1][36][86] = 1;dino_sprite[1][36][88] = 1;dino_sprite[1][36][89] = 1;dino_sprite[1][36][90] = 1;dino_sprite[1][36][91] = 1;dino_sprite[1][36][92] = 1;dino_sprite[1][37][44] = 1;dino_sprite[1][37][45] = 1;dino_sprite[1][37][46] = 1;dino_sprite[1][37][47] = 1;dino_sprite[1][37][48] = 1;dino_sprite[1][37][49] = 1;dino_sprite[1][37][50] = 1;dino_sprite[1][37][51] = 1;dino_sprite[1][37][52] = 1;dino_sprite[1][37][53] = 1;dino_sprite[1][37][54] = 1;dino_sprite[1][37][55] = 1;dino_sprite[1][37][56] = 1;dino_sprite[1][37][57] = 1;dino_sprite[1][37][58] = 1;dino_sprite[1][37][59] = 1;dino_sprite[1][37][60] = 1;dino_sprite[1][37][61] = 1;dino_sprite[1][37][62] = 1;dino_sprite[1][37][63] = 1;dino_sprite[1][37][64] = 1;dino_sprite[1][37][65] = 1;dino_sprite[1][37][66] = 1;dino_sprite[1][37][67] = 1;dino_sprite[1][37][68] = 1;dino_sprite[1][37][69] = 1;dino_sprite[1][37][70] = 1;dino_sprite[1][37][71] = 1;dino_sprite[1][37][72] = 1;dino_sprite[1][37][73] = 1;dino_sprite[1][37][74] = 1;dino_sprite[1][37][75] = 1;dino_sprite[1][37][76] = 1;dino_sprite[1][37][77] = 1;dino_sprite[1][37][78] = 1;dino_sprite[1][37][79] = 1;dino_sprite[1][37][80] = 1;dino_sprite[1][37][81] = 1;dino_sprite[1][37][82] = 1;dino_sprite[1][37][83] = 1;dino_sprite[1][37][84] = 1;dino_sprite[1][37][85] = 1;dino_sprite[1][37][86] = 1;dino_sprite[1][38][44] = 1;dino_sprite[1][38][45] = 1;dino_sprite[1][38][46] = 1;dino_sprite[1][38][47] = 1;dino_sprite[1][38][48] = 1;dino_sprite[1][38][49] = 1;dino_sprite[1][38][50] = 1;dino_sprite[1][38][51] = 1;dino_sprite[1][38][52] = 1;dino_sprite[1][38][53] = 1;dino_sprite[1][38][54] = 1;dino_sprite[1][38][55] = 1;dino_sprite[1][38][56] = 1;dino_sprite[1][38][57] = 1;dino_sprite[1][38][58] = 1;dino_sprite[1][38][59] = 1;dino_sprite[1][38][60] = 1;dino_sprite[1][38][61] = 1;dino_sprite[1][38][62] = 1;dino_sprite[1][38][63] = 1;dino_sprite[1][38][64] = 1;dino_sprite[1][38][65] = 1;dino_sprite[1][38][66] = 1;dino_sprite[1][38][67] = 1;dino_sprite[1][38][68] = 1;dino_sprite[1][38][69] = 1;dino_sprite[1][38][70] = 1;dino_sprite[1][38][71] = 1;dino_sprite[1][38][72] = 1;dino_sprite[1][38][73] = 1;dino_sprite[1][38][74] = 1;dino_sprite[1][38][75] = 1;dino_sprite[1][38][76] = 1;dino_sprite[1][38][77] = 1;dino_sprite[1][38][78] = 1;dino_sprite[1][38][79] = 1;dino_sprite[1][38][80] = 1;dino_sprite[1][38][81] = 1;dino_sprite[1][38][82] = 1;dino_sprite[1][38][83] = 1;dino_sprite[1][38][84] = 1;dino_sprite[1][38][85] = 1;dino_sprite[1][38][86] = 1;dino_sprite[1][39][39] = 1;dino_sprite[1][39][40] = 1;dino_sprite[1][39][41] = 1;dino_sprite[1][39][42] = 1;dino_sprite[1][39][43] = 1;dino_sprite[1][39][44] = 1;dino_sprite[1][39][45] = 1;dino_sprite[1][39][46] = 1;dino_sprite[1][39][47] = 1;dino_sprite[1][39][48] = 1;dino_sprite[1][39][49] = 1;dino_sprite[1][39][50] = 1;dino_sprite[1][39][51] = 1;dino_sprite[1][39][52] = 1;dino_sprite[1][39][53] = 1;dino_sprite[1][39][54] = 1;dino_sprite[1][39][55] = 1;dino_sprite[1][39][56] = 1;dino_sprite[1][39][57] = 1;dino_sprite[1][39][58] = 1;dino_sprite[1][39][59] = 1;dino_sprite[1][39][60] = 1;dino_sprite[1][39][61] = 1;dino_sprite[1][39][62] = 1;dino_sprite[1][39][63] = 1;dino_sprite[1][39][64] = 1;dino_sprite[1][39][65] = 1;dino_sprite[1][39][66] = 1;dino_sprite[1][39][67] = 1;dino_sprite[1][39][68] = 1;dino_sprite[1][39][69] = 1;dino_sprite[1][39][70] = 1;dino_sprite[1][39][71] = 1;dino_sprite[1][39][72] = 1;dino_sprite[1][39][73] = 1;dino_sprite[1][39][74] = 1;dino_sprite[1][39][75] = 1;dino_sprite[1][39][76] = 1;dino_sprite[1][39][77] = 1;dino_sprite[1][39][78] = 1;dino_sprite[1][39][79] = 1;dino_sprite[1][39][80] = 1;dino_sprite[1][39][81] = 1;dino_sprite[1][39][82] = 1;dino_sprite[1][39][83] = 1;dino_sprite[1][39][84] = 1;dino_sprite[1][39][85] = 1;dino_sprite[1][39][86] = 1;dino_sprite[1][40][39] = 1;dino_sprite[1][40][40] = 1;dino_sprite[1][40][41] = 1;dino_sprite[1][40][42] = 1;dino_sprite[1][40][43] = 1;dino_sprite[1][40][44] = 1;dino_sprite[1][40][45] = 1;dino_sprite[1][40][46] = 1;dino_sprite[1][40][47] = 1;dino_sprite[1][40][48] = 1;dino_sprite[1][40][49] = 1;dino_sprite[1][40][50] = 1;dino_sprite[1][40][51] = 1;dino_sprite[1][40][52] = 1;dino_sprite[1][40][53] = 1;dino_sprite[1][40][54] = 1;dino_sprite[1][40][55] = 1;dino_sprite[1][40][56] = 1;dino_sprite[1][40][57] = 1;dino_sprite[1][40][58] = 1;dino_sprite[1][40][59] = 1;dino_sprite[1][40][60] = 1;dino_sprite[1][40][61] = 1;dino_sprite[1][40][62] = 1;dino_sprite[1][40][63] = 1;dino_sprite[1][40][64] = 1;dino_sprite[1][40][65] = 1;dino_sprite[1][40][66] = 1;dino_sprite[1][40][67] = 1;dino_sprite[1][40][68] = 1;dino_sprite[1][40][69] = 1;dino_sprite[1][40][70] = 1;dino_sprite[1][40][71] = 1;dino_sprite[1][40][72] = 1;dino_sprite[1][40][73] = 1;dino_sprite[1][40][74] = 1;dino_sprite[1][40][75] = 1;dino_sprite[1][40][76] = 1;dino_sprite[1][40][77] = 1;dino_sprite[1][40][78] = 1;dino_sprite[1][40][79] = 1;dino_sprite[1][40][80] = 1;dino_sprite[1][40][81] = 1;dino_sprite[1][40][82] = 1;dino_sprite[1][40][83] = 1;dino_sprite[1][40][84] = 1;dino_sprite[1][40][85] = 1;dino_sprite[1][40][86] = 1;dino_sprite[1][41][39] = 1;dino_sprite[1][41][40] = 1;dino_sprite[1][41][41] = 1;dino_sprite[1][41][42] = 1;dino_sprite[1][41][43] = 1;dino_sprite[1][41][44] = 1;dino_sprite[1][41][45] = 1;dino_sprite[1][41][46] = 1;dino_sprite[1][41][47] = 1;dino_sprite[1][41][48] = 1;dino_sprite[1][41][49] = 1;dino_sprite[1][41][50] = 1;dino_sprite[1][41][51] = 1;dino_sprite[1][41][52] = 1;dino_sprite[1][41][53] = 1;dino_sprite[1][41][54] = 1;dino_sprite[1][41][55] = 1;dino_sprite[1][41][56] = 1;dino_sprite[1][41][57] = 1;dino_sprite[1][41][58] = 1;dino_sprite[1][41][59] = 1;dino_sprite[1][41][60] = 1;dino_sprite[1][41][61] = 1;dino_sprite[1][41][62] = 1;dino_sprite[1][41][63] = 1;dino_sprite[1][41][64] = 1;dino_sprite[1][41][65] = 1;dino_sprite[1][41][66] = 1;dino_sprite[1][41][67] = 1;dino_sprite[1][41][68] = 1;dino_sprite[1][41][69] = 1;dino_sprite[1][41][70] = 1;dino_sprite[1][41][71] = 1;dino_sprite[1][41][72] = 1;dino_sprite[1][41][73] = 1;dino_sprite[1][41][74] = 1;dino_sprite[1][41][75] = 1;dino_sprite[1][41][76] = 1;dino_sprite[1][41][77] = 1;dino_sprite[1][41][78] = 1;dino_sprite[1][41][79] = 1;dino_sprite[1][41][80] = 1;dino_sprite[1][41][81] = 1;dino_sprite[1][41][82] = 1;dino_sprite[1][42][39] = 1;dino_sprite[1][42][40] = 1;dino_sprite[1][42][41] = 1;dino_sprite[1][42][42] = 1;dino_sprite[1][42][43] = 1;dino_sprite[1][42][44] = 1;dino_sprite[1][42][45] = 1;dino_sprite[1][42][46] = 1;dino_sprite[1][42][47] = 1;dino_sprite[1][42][48] = 1;dino_sprite[1][42][49] = 1;dino_sprite[1][42][50] = 1;dino_sprite[1][42][51] = 1;dino_sprite[1][42][52] = 1;dino_sprite[1][42][53] = 1;dino_sprite[1][42][54] = 1;dino_sprite[1][42][55] = 1;dino_sprite[1][42][56] = 1;dino_sprite[1][42][57] = 1;dino_sprite[1][42][58] = 1;dino_sprite[1][42][59] = 1;dino_sprite[1][42][60] = 1;dino_sprite[1][42][61] = 1;dino_sprite[1][42][62] = 1;dino_sprite[1][42][63] = 1;dino_sprite[1][42][64] = 1;dino_sprite[1][42][65] = 1;dino_sprite[1][42][66] = 1;dino_sprite[1][42][67] = 1;dino_sprite[1][42][68] = 1;dino_sprite[1][42][69] = 1;dino_sprite[1][42][70] = 1;dino_sprite[1][42][71] = 1;dino_sprite[1][42][72] = 1;dino_sprite[1][42][73] = 1;dino_sprite[1][42][74] = 1;dino_sprite[1][42][75] = 1;dino_sprite[1][42][76] = 1;dino_sprite[1][42][77] = 1;dino_sprite[1][42][78] = 1;dino_sprite[1][42][79] = 1;dino_sprite[1][42][80] = 1;dino_sprite[1][42][81] = 1;dino_sprite[1][42][82] = 1;dino_sprite[1][43][39] = 1;dino_sprite[1][43][40] = 1;dino_sprite[1][43][41] = 1;dino_sprite[1][43][42] = 1;dino_sprite[1][43][43] = 1;dino_sprite[1][43][44] = 1;dino_sprite[1][43][45] = 1;dino_sprite[1][43][46] = 1;dino_sprite[1][43][47] = 1;dino_sprite[1][43][48] = 1;dino_sprite[1][43][49] = 1;dino_sprite[1][43][50] = 1;dino_sprite[1][43][51] = 1;dino_sprite[1][43][52] = 1;dino_sprite[1][43][53] = 1;dino_sprite[1][43][54] = 1;dino_sprite[1][43][55] = 1;dino_sprite[1][43][56] = 1;dino_sprite[1][43][57] = 1;dino_sprite[1][43][58] = 1;dino_sprite[1][43][59] = 1;dino_sprite[1][43][60] = 1;dino_sprite[1][43][61] = 1;dino_sprite[1][43][62] = 1;dino_sprite[1][43][63] = 1;dino_sprite[1][43][64] = 1;dino_sprite[1][43][65] = 1;dino_sprite[1][43][66] = 1;dino_sprite[1][43][67] = 1;dino_sprite[1][43][68] = 1;dino_sprite[1][43][69] = 1;dino_sprite[1][43][70] = 1;dino_sprite[1][43][71] = 1;dino_sprite[1][43][72] = 1;dino_sprite[1][43][73] = 1;dino_sprite[1][43][74] = 1;dino_sprite[1][43][75] = 1;dino_sprite[1][43][76] = 1;dino_sprite[1][43][77] = 1;dino_sprite[1][43][78] = 1;dino_sprite[1][43][79] = 1;dino_sprite[1][43][80] = 1;dino_sprite[1][43][81] = 1;dino_sprite[1][43][82] = 1;dino_sprite[1][44][39] = 1;dino_sprite[1][44][40] = 1;dino_sprite[1][44][41] = 1;dino_sprite[1][44][42] = 1;dino_sprite[1][44][43] = 1;dino_sprite[1][44][44] = 1;dino_sprite[1][44][45] = 1;dino_sprite[1][44][46] = 1;dino_sprite[1][44][47] = 1;dino_sprite[1][44][48] = 1;dino_sprite[1][44][49] = 1;dino_sprite[1][44][50] = 1;dino_sprite[1][44][51] = 1;dino_sprite[1][44][52] = 1;dino_sprite[1][44][53] = 1;dino_sprite[1][44][54] = 1;dino_sprite[1][44][55] = 1;dino_sprite[1][44][56] = 1;dino_sprite[1][44][57] = 1;dino_sprite[1][44][58] = 1;dino_sprite[1][44][59] = 1;dino_sprite[1][44][60] = 1;dino_sprite[1][44][61] = 1;dino_sprite[1][44][62] = 1;dino_sprite[1][44][63] = 1;dino_sprite[1][44][64] = 1;dino_sprite[1][44][65] = 1;dino_sprite[1][44][66] = 1;dino_sprite[1][44][67] = 1;dino_sprite[1][44][68] = 1;dino_sprite[1][44][69] = 1;dino_sprite[1][44][70] = 1;dino_sprite[1][44][71] = 1;dino_sprite[1][44][72] = 1;dino_sprite[1][44][73] = 1;dino_sprite[1][44][74] = 1;dino_sprite[1][44][75] = 1;dino_sprite[1][44][76] = 1;dino_sprite[1][44][77] = 1;dino_sprite[1][44][78] = 1;dino_sprite[1][44][79] = 1;dino_sprite[1][44][80] = 1;dino_sprite[1][44][81] = 1;dino_sprite[1][44][82] = 1;dino_sprite[1][45][35] = 1;dino_sprite[1][45][36] = 1;dino_sprite[1][45][37] = 1;dino_sprite[1][45][39] = 1;dino_sprite[1][45][40] = 1;dino_sprite[1][45][41] = 1;dino_sprite[1][45][42] = 1;dino_sprite[1][45][43] = 1;dino_sprite[1][45][44] = 1;dino_sprite[1][45][45] = 1;dino_sprite[1][45][46] = 1;dino_sprite[1][45][47] = 1;dino_sprite[1][45][48] = 1;dino_sprite[1][45][49] = 1;dino_sprite[1][45][50] = 1;dino_sprite[1][45][51] = 1;dino_sprite[1][45][52] = 1;dino_sprite[1][45][53] = 1;dino_sprite[1][45][54] = 1;dino_sprite[1][45][55] = 1;dino_sprite[1][45][56] = 1;dino_sprite[1][45][57] = 1;dino_sprite[1][45][58] = 1;dino_sprite[1][45][59] = 1;dino_sprite[1][45][60] = 1;dino_sprite[1][45][61] = 1;dino_sprite[1][45][62] = 1;dino_sprite[1][45][63] = 1;dino_sprite[1][45][64] = 1;dino_sprite[1][45][65] = 1;dino_sprite[1][45][66] = 1;dino_sprite[1][45][67] = 1;dino_sprite[1][45][68] = 1;dino_sprite[1][45][69] = 1;dino_sprite[1][45][70] = 1;dino_sprite[1][45][71] = 1;dino_sprite[1][45][72] = 1;dino_sprite[1][45][73] = 1;dino_sprite[1][45][74] = 1;dino_sprite[1][45][75] = 1;dino_sprite[1][45][76] = 1;dino_sprite[1][45][77] = 1;dino_sprite[1][45][78] = 1;dino_sprite[1][45][79] = 1;dino_sprite[1][45][80] = 1;dino_sprite[1][45][81] = 1;dino_sprite[1][45][82] = 1;dino_sprite[1][45][84] = 1;dino_sprite[1][45][85] = 1;dino_sprite[1][45][86] = 1;dino_sprite[1][46][35] = 1;dino_sprite[1][46][36] = 1;dino_sprite[1][46][37] = 1;dino_sprite[1][46][38] = 1;dino_sprite[1][46][39] = 1;dino_sprite[1][46][40] = 1;dino_sprite[1][46][41] = 1;dino_sprite[1][46][42] = 1;dino_sprite[1][46][43] = 1;dino_sprite[1][46][44] = 1;dino_sprite[1][46][45] = 1;dino_sprite[1][46][46] = 1;dino_sprite[1][46][47] = 1;dino_sprite[1][46][48] = 1;dino_sprite[1][46][49] = 1;dino_sprite[1][46][50] = 1;dino_sprite[1][46][51] = 1;dino_sprite[1][46][52] = 1;dino_sprite[1][46][53] = 1;dino_sprite[1][46][54] = 1;dino_sprite[1][46][55] = 1;dino_sprite[1][46][56] = 1;dino_sprite[1][46][57] = 1;dino_sprite[1][46][58] = 1;dino_sprite[1][46][59] = 1;dino_sprite[1][46][60] = 1;dino_sprite[1][46][61] = 1;dino_sprite[1][46][62] = 1;dino_sprite[1][46][63] = 1;dino_sprite[1][46][64] = 1;dino_sprite[1][46][65] = 1;dino_sprite[1][46][66] = 1;dino_sprite[1][46][67] = 1;dino_sprite[1][46][68] = 1;dino_sprite[1][46][69] = 1;dino_sprite[1][46][70] = 1;dino_sprite[1][46][71] = 1;dino_sprite[1][46][72] = 1;dino_sprite[1][46][73] = 1;dino_sprite[1][46][74] = 1;dino_sprite[1][46][75] = 1;dino_sprite[1][46][76] = 1;dino_sprite[1][46][77] = 1;dino_sprite[1][46][78] = 1;dino_sprite[1][46][79] = 1;dino_sprite[1][46][80] = 1;dino_sprite[1][46][81] = 1;dino_sprite[1][46][82] = 1;dino_sprite[1][46][83] = 1;dino_sprite[1][46][84] = 1;dino_sprite[1][46][85] = 1;dino_sprite[1][46][86] = 1;dino_sprite[1][47][35] = 1;dino_sprite[1][47][36] = 1;dino_sprite[1][47][37] = 1;dino_sprite[1][47][38] = 1;dino_sprite[1][47][39] = 1;dino_sprite[1][47][40] = 1;dino_sprite[1][47][41] = 1;dino_sprite[1][47][42] = 1;dino_sprite[1][47][43] = 1;dino_sprite[1][47][44] = 1;dino_sprite[1][47][45] = 1;dino_sprite[1][47][46] = 1;dino_sprite[1][47][47] = 1;dino_sprite[1][47][48] = 1;dino_sprite[1][47][49] = 1;dino_sprite[1][47][50] = 1;dino_sprite[1][47][51] = 1;dino_sprite[1][47][52] = 1;dino_sprite[1][47][53] = 1;dino_sprite[1][47][54] = 1;dino_sprite[1][47][55] = 1;dino_sprite[1][47][56] = 1;dino_sprite[1][47][57] = 1;dino_sprite[1][47][58] = 1;dino_sprite[1][47][59] = 1;dino_sprite[1][47][60] = 1;dino_sprite[1][47][61] = 1;dino_sprite[1][47][62] = 1;dino_sprite[1][47][63] = 1;dino_sprite[1][47][64] = 1;dino_sprite[1][47][65] = 1;dino_sprite[1][47][66] = 1;dino_sprite[1][47][67] = 1;dino_sprite[1][47][68] = 1;dino_sprite[1][47][69] = 1;dino_sprite[1][47][70] = 1;dino_sprite[1][47][71] = 1;dino_sprite[1][47][72] = 1;dino_sprite[1][47][73] = 1;dino_sprite[1][47][74] = 1;dino_sprite[1][47][75] = 1;dino_sprite[1][47][76] = 1;dino_sprite[1][47][77] = 1;dino_sprite[1][47][78] = 1;dino_sprite[1][47][79] = 1;dino_sprite[1][47][80] = 1;dino_sprite[1][47][81] = 1;dino_sprite[1][47][82] = 1;dino_sprite[1][47][83] = 1;dino_sprite[1][47][84] = 1;dino_sprite[1][47][85] = 1;dino_sprite[1][47][86] = 1;dino_sprite[1][48][35] = 1;dino_sprite[1][48][36] = 1;dino_sprite[1][48][37] = 1;dino_sprite[1][48][38] = 1;dino_sprite[1][48][39] = 1;dino_sprite[1][48][40] = 1;dino_sprite[1][48][41] = 1;dino_sprite[1][48][42] = 1;dino_sprite[1][48][43] = 1;dino_sprite[1][48][44] = 1;dino_sprite[1][48][45] = 1;dino_sprite[1][48][46] = 1;dino_sprite[1][48][47] = 1;dino_sprite[1][48][48] = 1;dino_sprite[1][48][49] = 1;dino_sprite[1][48][50] = 1;dino_sprite[1][48][51] = 1;dino_sprite[1][48][52] = 1;dino_sprite[1][48][53] = 1;dino_sprite[1][48][54] = 1;dino_sprite[1][48][55] = 1;dino_sprite[1][48][56] = 1;dino_sprite[1][48][57] = 1;dino_sprite[1][48][58] = 1;dino_sprite[1][48][59] = 1;dino_sprite[1][48][60] = 1;dino_sprite[1][48][61] = 1;dino_sprite[1][48][62] = 1;dino_sprite[1][48][63] = 1;dino_sprite[1][48][64] = 1;dino_sprite[1][48][65] = 1;dino_sprite[1][48][66] = 1;dino_sprite[1][48][67] = 1;dino_sprite[1][48][68] = 1;dino_sprite[1][48][69] = 1;dino_sprite[1][48][70] = 1;dino_sprite[1][48][71] = 1;dino_sprite[1][48][72] = 1;dino_sprite[1][48][73] = 1;dino_sprite[1][48][74] = 1;dino_sprite[1][48][75] = 1;dino_sprite[1][48][76] = 1;dino_sprite[1][48][77] = 1;dino_sprite[1][48][78] = 1;dino_sprite[1][48][79] = 1;dino_sprite[1][48][80] = 1;dino_sprite[1][48][81] = 1;dino_sprite[1][48][82] = 1;dino_sprite[1][48][83] = 1;dino_sprite[1][48][84] = 1;dino_sprite[1][48][85] = 1;dino_sprite[1][48][86] = 1;dino_sprite[1][49][35] = 1;dino_sprite[1][49][36] = 1;dino_sprite[1][49][37] = 1;dino_sprite[1][49][38] = 1;dino_sprite[1][49][39] = 1;dino_sprite[1][49][40] = 1;dino_sprite[1][49][41] = 1;dino_sprite[1][49][42] = 1;dino_sprite[1][49][43] = 1;dino_sprite[1][49][44] = 1;dino_sprite[1][49][45] = 1;dino_sprite[1][49][46] = 1;dino_sprite[1][49][47] = 1;dino_sprite[1][49][48] = 1;dino_sprite[1][49][49] = 1;dino_sprite[1][49][50] = 1;dino_sprite[1][49][51] = 1;dino_sprite[1][49][52] = 1;dino_sprite[1][49][53] = 1;dino_sprite[1][49][54] = 1;dino_sprite[1][49][55] = 1;dino_sprite[1][49][56] = 1;dino_sprite[1][49][57] = 1;dino_sprite[1][49][58] = 1;dino_sprite[1][49][59] = 1;dino_sprite[1][49][60] = 1;dino_sprite[1][49][61] = 1;dino_sprite[1][49][62] = 1;dino_sprite[1][49][63] = 1;dino_sprite[1][49][64] = 1;dino_sprite[1][49][65] = 1;dino_sprite[1][49][66] = 1;dino_sprite[1][49][67] = 1;dino_sprite[1][49][68] = 1;dino_sprite[1][49][69] = 1;dino_sprite[1][49][70] = 1;dino_sprite[1][49][71] = 1;dino_sprite[1][49][72] = 1;dino_sprite[1][49][73] = 1;dino_sprite[1][49][74] = 1;dino_sprite[1][49][75] = 1;dino_sprite[1][49][76] = 1;dino_sprite[1][49][77] = 1;dino_sprite[1][49][78] = 1;dino_sprite[1][49][79] = 1;dino_sprite[1][49][80] = 1;dino_sprite[1][49][81] = 1;dino_sprite[1][49][82] = 1;dino_sprite[1][49][83] = 1;dino_sprite[1][49][84] = 1;dino_sprite[1][49][85] = 1;dino_sprite[1][49][86] = 1;dino_sprite[1][50][35] = 1;dino_sprite[1][50][36] = 1;dino_sprite[1][50][37] = 1;dino_sprite[1][50][38] = 1;dino_sprite[1][50][39] = 1;dino_sprite[1][50][40] = 1;dino_sprite[1][50][41] = 1;dino_sprite[1][50][42] = 1;dino_sprite[1][50][43] = 1;dino_sprite[1][50][44] = 1;dino_sprite[1][50][45] = 1;dino_sprite[1][50][46] = 1;dino_sprite[1][50][47] = 1;dino_sprite[1][50][48] = 1;dino_sprite[1][50][49] = 1;dino_sprite[1][50][50] = 1;dino_sprite[1][50][51] = 1;dino_sprite[1][50][52] = 1;dino_sprite[1][50][53] = 1;dino_sprite[1][50][54] = 1;dino_sprite[1][50][55] = 1;dino_sprite[1][50][56] = 1;dino_sprite[1][50][57] = 1;dino_sprite[1][50][58] = 1;dino_sprite[1][50][59] = 1;dino_sprite[1][50][60] = 1;dino_sprite[1][50][61] = 1;dino_sprite[1][50][62] = 1;dino_sprite[1][50][63] = 1;dino_sprite[1][50][64] = 1;dino_sprite[1][50][65] = 1;dino_sprite[1][50][66] = 1;dino_sprite[1][50][67] = 1;dino_sprite[1][50][68] = 1;dino_sprite[1][50][69] = 1;dino_sprite[1][50][70] = 1;dino_sprite[1][50][71] = 1;dino_sprite[1][50][72] = 1;dino_sprite[1][50][73] = 1;dino_sprite[1][50][74] = 1;dino_sprite[1][50][75] = 1;dino_sprite[1][50][76] = 1;dino_sprite[1][50][77] = 1;dino_sprite[1][50][78] = 1;dino_sprite[1][50][79] = 1;dino_sprite[1][50][80] = 1;dino_sprite[1][50][81] = 1;dino_sprite[1][50][82] = 1;dino_sprite[1][50][83] = 1;dino_sprite[1][50][84] = 1;dino_sprite[1][50][85] = 1;dino_sprite[1][50][86] = 1;dino_sprite[1][50][88] = 1;dino_sprite[1][50][89] = 1;dino_sprite[1][50][90] = 1;dino_sprite[1][50][91] = 1;dino_sprite[1][50][92] = 1;dino_sprite[1][50][93] = 1;dino_sprite[1][50][94] = 1;dino_sprite[1][50][95] = 1;dino_sprite[1][50][96] = 1;dino_sprite[1][50][97] = 1;dino_sprite[1][50][98] = 1;dino_sprite[1][50][99] = 1;dino_sprite[1][51][3] = 1;dino_sprite[1][51][4] = 1;dino_sprite[1][51][5] = 1;dino_sprite[1][51][6] = 1;dino_sprite[1][51][7] = 1;dino_sprite[1][51][8] = 1;dino_sprite[1][51][9] = 1;dino_sprite[1][51][10] = 1;dino_sprite[1][51][11] = 1;dino_sprite[1][51][12] = 1;dino_sprite[1][51][13] = 1;dino_sprite[1][51][14] = 1;dino_sprite[1][51][15] = 1;dino_sprite[1][51][16] = 1;dino_sprite[1][51][17] = 1;dino_sprite[1][51][18] = 1;dino_sprite[1][51][19] = 1;dino_sprite[1][51][20] = 1;dino_sprite[1][51][21] = 1;dino_sprite[1][51][22] = 1;dino_sprite[1][51][23] = 1;dino_sprite[1][51][24] = 1;dino_sprite[1][51][25] = 1;dino_sprite[1][51][26] = 1;dino_sprite[1][51][27] = 1;dino_sprite[1][51][28] = 1;dino_sprite[1][51][29] = 1;dino_sprite[1][51][30] = 1;dino_sprite[1][51][31] = 1;dino_sprite[1][51][32] = 1;dino_sprite[1][51][33] = 1;dino_sprite[1][51][34] = 1;dino_sprite[1][51][35] = 1;dino_sprite[1][51][36] = 1;dino_sprite[1][51][37] = 1;dino_sprite[1][51][38] = 1;dino_sprite[1][51][39] = 1;dino_sprite[1][51][40] = 1;dino_sprite[1][51][41] = 1;dino_sprite[1][51][42] = 1;dino_sprite[1][51][43] = 1;dino_sprite[1][51][44] = 1;dino_sprite[1][51][45] = 1;dino_sprite[1][51][46] = 1;dino_sprite[1][51][47] = 1;dino_sprite[1][51][48] = 1;dino_sprite[1][51][49] = 1;dino_sprite[1][51][50] = 1;dino_sprite[1][51][51] = 1;dino_sprite[1][51][52] = 1;dino_sprite[1][51][53] = 1;dino_sprite[1][51][54] = 1;dino_sprite[1][51][55] = 1;dino_sprite[1][51][56] = 1;dino_sprite[1][51][57] = 1;dino_sprite[1][51][58] = 1;dino_sprite[1][51][59] = 1;dino_sprite[1][51][60] = 1;dino_sprite[1][51][61] = 1;dino_sprite[1][51][62] = 1;dino_sprite[1][51][63] = 1;dino_sprite[1][51][64] = 1;dino_sprite[1][51][65] = 1;dino_sprite[1][51][66] = 1;dino_sprite[1][51][67] = 1;dino_sprite[1][51][68] = 1;dino_sprite[1][51][69] = 1;dino_sprite[1][51][70] = 1;dino_sprite[1][51][71] = 1;dino_sprite[1][51][72] = 1;dino_sprite[1][51][73] = 1;dino_sprite[1][51][74] = 1;dino_sprite[1][51][75] = 1;dino_sprite[1][51][76] = 1;dino_sprite[1][51][77] = 1;dino_sprite[1][51][78] = 1;dino_sprite[1][51][79] = 1;dino_sprite[1][51][80] = 1;dino_sprite[1][51][81] = 1;dino_sprite[1][51][82] = 1;dino_sprite[1][51][83] = 1;dino_sprite[1][51][84] = 1;dino_sprite[1][51][85] = 1;dino_sprite[1][51][86] = 1;dino_sprite[1][51][87] = 1;dino_sprite[1][51][88] = 1;dino_sprite[1][51][89] = 1;dino_sprite[1][51][90] = 1;dino_sprite[1][51][91] = 1;dino_sprite[1][51][92] = 1;dino_sprite[1][51][93] = 1;dino_sprite[1][51][94] = 1;dino_sprite[1][51][95] = 1;dino_sprite[1][51][96] = 1;dino_sprite[1][51][97] = 1;dino_sprite[1][51][98] = 1;dino_sprite[1][51][99] = 1;dino_sprite[1][52][3] = 1;dino_sprite[1][52][4] = 1;dino_sprite[1][52][5] = 1;dino_sprite[1][52][6] = 1;dino_sprite[1][52][7] = 1;dino_sprite[1][52][8] = 1;dino_sprite[1][52][9] = 1;dino_sprite[1][52][10] = 1;dino_sprite[1][52][11] = 1;dino_sprite[1][52][12] = 1;dino_sprite[1][52][13] = 1;dino_sprite[1][52][14] = 1;dino_sprite[1][52][15] = 1;dino_sprite[1][52][16] = 1;dino_sprite[1][52][17] = 1;dino_sprite[1][52][18] = 1;dino_sprite[1][52][19] = 1;dino_sprite[1][52][20] = 1;dino_sprite[1][52][21] = 1;dino_sprite[1][52][22] = 1;dino_sprite[1][52][23] = 1;dino_sprite[1][52][24] = 1;dino_sprite[1][52][25] = 1;dino_sprite[1][52][26] = 1;dino_sprite[1][52][27] = 1;dino_sprite[1][52][28] = 1;dino_sprite[1][52][29] = 1;dino_sprite[1][52][30] = 1;dino_sprite[1][52][31] = 1;dino_sprite[1][52][32] = 1;dino_sprite[1][52][33] = 1;dino_sprite[1][52][34] = 1;dino_sprite[1][52][35] = 1;dino_sprite[1][52][36] = 1;dino_sprite[1][52][37] = 1;dino_sprite[1][52][38] = 1;dino_sprite[1][52][39] = 1;dino_sprite[1][52][40] = 1;dino_sprite[1][52][41] = 1;dino_sprite[1][52][42] = 1;dino_sprite[1][52][43] = 1;dino_sprite[1][52][44] = 1;dino_sprite[1][52][45] = 1;dino_sprite[1][52][46] = 1;dino_sprite[1][52][47] = 1;dino_sprite[1][52][48] = 1;dino_sprite[1][52][49] = 1;dino_sprite[1][52][50] = 1;dino_sprite[1][52][51] = 1;dino_sprite[1][52][52] = 1;dino_sprite[1][52][53] = 1;dino_sprite[1][52][54] = 1;dino_sprite[1][52][55] = 1;dino_sprite[1][52][56] = 1;dino_sprite[1][52][57] = 1;dino_sprite[1][52][58] = 1;dino_sprite[1][52][59] = 1;dino_sprite[1][52][60] = 1;dino_sprite[1][52][61] = 1;dino_sprite[1][52][62] = 1;dino_sprite[1][52][63] = 1;dino_sprite[1][52][64] = 1;dino_sprite[1][52][65] = 1;dino_sprite[1][52][66] = 1;dino_sprite[1][52][67] = 1;dino_sprite[1][52][68] = 1;dino_sprite[1][52][69] = 1;dino_sprite[1][52][70] = 1;dino_sprite[1][52][71] = 1;dino_sprite[1][52][72] = 1;dino_sprite[1][52][73] = 1;dino_sprite[1][52][74] = 1;dino_sprite[1][52][75] = 1;dino_sprite[1][52][76] = 1;dino_sprite[1][52][77] = 1;dino_sprite[1][52][78] = 1;dino_sprite[1][52][79] = 1;dino_sprite[1][52][80] = 1;dino_sprite[1][52][81] = 1;dino_sprite[1][52][82] = 1;dino_sprite[1][52][83] = 1;dino_sprite[1][52][84] = 1;dino_sprite[1][52][85] = 1;dino_sprite[1][52][86] = 1;dino_sprite[1][52][87] = 1;dino_sprite[1][52][88] = 1;dino_sprite[1][52][89] = 1;dino_sprite[1][52][90] = 1;dino_sprite[1][52][91] = 1;dino_sprite[1][52][92] = 1;dino_sprite[1][52][93] = 1;dino_sprite[1][52][94] = 1;dino_sprite[1][52][95] = 1;dino_sprite[1][52][96] = 1;dino_sprite[1][52][97] = 1;dino_sprite[1][52][98] = 1;dino_sprite[1][52][99] = 1;dino_sprite[1][53][3] = 1;dino_sprite[1][53][4] = 1;dino_sprite[1][53][5] = 1;dino_sprite[1][53][6] = 1;dino_sprite[1][53][7] = 1;dino_sprite[1][53][8] = 1;dino_sprite[1][53][9] = 1;dino_sprite[1][53][10] = 1;dino_sprite[1][53][11] = 1;dino_sprite[1][53][12] = 1;dino_sprite[1][53][13] = 1;dino_sprite[1][53][14] = 1;dino_sprite[1][53][15] = 1;dino_sprite[1][53][16] = 1;dino_sprite[1][53][17] = 1;dino_sprite[1][53][18] = 1;dino_sprite[1][53][19] = 1;dino_sprite[1][53][20] = 1;dino_sprite[1][53][21] = 1;dino_sprite[1][53][22] = 1;dino_sprite[1][53][23] = 1;dino_sprite[1][53][24] = 1;dino_sprite[1][53][25] = 1;dino_sprite[1][53][26] = 1;dino_sprite[1][53][27] = 1;dino_sprite[1][53][28] = 1;dino_sprite[1][53][29] = 1;dino_sprite[1][53][30] = 1;dino_sprite[1][53][31] = 1;dino_sprite[1][53][32] = 1;dino_sprite[1][53][33] = 1;dino_sprite[1][53][34] = 1;dino_sprite[1][53][35] = 1;dino_sprite[1][53][36] = 1;dino_sprite[1][53][37] = 1;dino_sprite[1][53][38] = 1;dino_sprite[1][53][39] = 1;dino_sprite[1][53][40] = 1;dino_sprite[1][53][41] = 1;dino_sprite[1][53][42] = 1;dino_sprite[1][53][43] = 1;dino_sprite[1][53][44] = 1;dino_sprite[1][53][45] = 1;dino_sprite[1][53][46] = 1;dino_sprite[1][53][47] = 1;dino_sprite[1][53][48] = 1;dino_sprite[1][53][49] = 1;dino_sprite[1][53][50] = 1;dino_sprite[1][53][51] = 1;dino_sprite[1][53][52] = 1;dino_sprite[1][53][53] = 1;dino_sprite[1][53][54] = 1;dino_sprite[1][53][55] = 1;dino_sprite[1][53][56] = 1;dino_sprite[1][53][57] = 1;dino_sprite[1][53][58] = 1;dino_sprite[1][53][59] = 1;dino_sprite[1][53][60] = 1;dino_sprite[1][53][61] = 1;dino_sprite[1][53][62] = 1;dino_sprite[1][53][63] = 1;dino_sprite[1][53][64] = 1;dino_sprite[1][53][65] = 1;dino_sprite[1][53][66] = 1;dino_sprite[1][53][67] = 1;dino_sprite[1][53][68] = 1;dino_sprite[1][53][69] = 1;dino_sprite[1][53][70] = 1;dino_sprite[1][53][71] = 1;dino_sprite[1][53][72] = 1;dino_sprite[1][53][73] = 1;dino_sprite[1][53][74] = 1;dino_sprite[1][53][75] = 1;dino_sprite[1][53][76] = 1;dino_sprite[1][53][77] = 1;dino_sprite[1][53][78] = 1;dino_sprite[1][53][79] = 1;dino_sprite[1][53][80] = 1;dino_sprite[1][53][81] = 1;dino_sprite[1][53][82] = 1;dino_sprite[1][53][83] = 1;dino_sprite[1][53][84] = 1;dino_sprite[1][53][85] = 1;dino_sprite[1][53][86] = 1;dino_sprite[1][53][87] = 1;dino_sprite[1][53][88] = 1;dino_sprite[1][53][89] = 1;dino_sprite[1][53][90] = 1;dino_sprite[1][53][91] = 1;dino_sprite[1][53][92] = 1;dino_sprite[1][53][93] = 1;dino_sprite[1][53][94] = 1;dino_sprite[1][53][95] = 1;dino_sprite[1][53][96] = 1;dino_sprite[1][53][97] = 1;dino_sprite[1][53][98] = 1;dino_sprite[1][53][99] = 1;dino_sprite[1][54][3] = 1;dino_sprite[1][54][4] = 1;dino_sprite[1][54][5] = 1;dino_sprite[1][54][6] = 1;dino_sprite[1][54][7] = 1;dino_sprite[1][54][8] = 1;dino_sprite[1][54][9] = 1;dino_sprite[1][54][10] = 1;dino_sprite[1][54][11] = 1;dino_sprite[1][54][12] = 1;dino_sprite[1][54][13] = 1;dino_sprite[1][54][14] = 1;dino_sprite[1][54][15] = 1;dino_sprite[1][54][16] = 1;dino_sprite[1][54][17] = 1;dino_sprite[1][54][18] = 1;dino_sprite[1][54][19] = 1;dino_sprite[1][54][20] = 1;dino_sprite[1][54][21] = 1;dino_sprite[1][54][22] = 1;dino_sprite[1][54][23] = 1;dino_sprite[1][54][24] = 1;dino_sprite[1][54][25] = 1;dino_sprite[1][54][26] = 1;dino_sprite[1][54][27] = 1;dino_sprite[1][54][28] = 1;dino_sprite[1][54][29] = 1;dino_sprite[1][54][30] = 1;dino_sprite[1][54][31] = 1;dino_sprite[1][54][32] = 1;dino_sprite[1][54][33] = 1;dino_sprite[1][54][34] = 1;dino_sprite[1][54][35] = 1;dino_sprite[1][54][36] = 1;dino_sprite[1][54][37] = 1;dino_sprite[1][54][38] = 1;dino_sprite[1][54][39] = 1;dino_sprite[1][54][40] = 1;dino_sprite[1][54][41] = 1;dino_sprite[1][54][42] = 1;dino_sprite[1][54][43] = 1;dino_sprite[1][54][44] = 1;dino_sprite[1][54][45] = 1;dino_sprite[1][54][46] = 1;dino_sprite[1][54][47] = 1;dino_sprite[1][54][48] = 1;dino_sprite[1][54][49] = 1;dino_sprite[1][54][50] = 1;dino_sprite[1][54][51] = 1;dino_sprite[1][54][52] = 1;dino_sprite[1][54][53] = 1;dino_sprite[1][54][54] = 1;dino_sprite[1][54][55] = 1;dino_sprite[1][54][56] = 1;dino_sprite[1][54][57] = 1;dino_sprite[1][54][58] = 1;dino_sprite[1][54][59] = 1;dino_sprite[1][54][60] = 1;dino_sprite[1][54][61] = 1;dino_sprite[1][54][62] = 1;dino_sprite[1][54][63] = 1;dino_sprite[1][54][64] = 1;dino_sprite[1][54][65] = 1;dino_sprite[1][54][66] = 1;dino_sprite[1][54][67] = 1;dino_sprite[1][54][68] = 1;dino_sprite[1][54][69] = 1;dino_sprite[1][54][70] = 1;dino_sprite[1][54][71] = 1;dino_sprite[1][54][72] = 1;dino_sprite[1][54][73] = 1;dino_sprite[1][54][74] = 1;dino_sprite[1][54][75] = 1;dino_sprite[1][54][76] = 1;dino_sprite[1][54][77] = 1;dino_sprite[1][54][78] = 1;dino_sprite[1][54][79] = 1;dino_sprite[1][54][80] = 1;dino_sprite[1][54][81] = 1;dino_sprite[1][54][82] = 1;dino_sprite[1][54][83] = 1;dino_sprite[1][54][84] = 1;dino_sprite[1][54][85] = 1;dino_sprite[1][54][86] = 1;dino_sprite[1][54][87] = 1;dino_sprite[1][54][88] = 1;dino_sprite[1][54][89] = 1;dino_sprite[1][54][90] = 1;dino_sprite[1][54][91] = 1;dino_sprite[1][54][92] = 1;dino_sprite[1][54][93] = 1;dino_sprite[1][54][94] = 1;dino_sprite[1][54][95] = 1;dino_sprite[1][54][96] = 1;dino_sprite[1][54][97] = 1;dino_sprite[1][54][98] = 1;dino_sprite[1][54][99] = 1;dino_sprite[1][55][3] = 1;dino_sprite[1][55][4] = 1;dino_sprite[1][55][5] = 1;dino_sprite[1][55][6] = 1;dino_sprite[1][55][7] = 1;dino_sprite[1][55][8] = 1;dino_sprite[1][55][9] = 1;dino_sprite[1][55][10] = 1;dino_sprite[1][55][11] = 1;dino_sprite[1][55][12] = 1;dino_sprite[1][55][13] = 1;dino_sprite[1][55][14] = 1;dino_sprite[1][55][15] = 1;dino_sprite[1][55][16] = 1;dino_sprite[1][55][17] = 1;dino_sprite[1][55][18] = 1;dino_sprite[1][55][19] = 1;dino_sprite[1][55][20] = 1;dino_sprite[1][55][21] = 1;dino_sprite[1][55][22] = 1;dino_sprite[1][55][23] = 1;dino_sprite[1][55][24] = 1;dino_sprite[1][55][25] = 1;dino_sprite[1][55][26] = 1;dino_sprite[1][55][27] = 1;dino_sprite[1][55][28] = 1;dino_sprite[1][55][29] = 1;dino_sprite[1][55][30] = 1;dino_sprite[1][55][31] = 1;dino_sprite[1][55][32] = 1;dino_sprite[1][55][33] = 1;dino_sprite[1][55][34] = 1;dino_sprite[1][55][35] = 1;dino_sprite[1][55][36] = 1;dino_sprite[1][55][37] = 1;dino_sprite[1][55][38] = 1;dino_sprite[1][55][39] = 1;dino_sprite[1][55][40] = 1;dino_sprite[1][55][41] = 1;dino_sprite[1][55][42] = 1;dino_sprite[1][55][43] = 1;dino_sprite[1][55][44] = 1;dino_sprite[1][55][45] = 1;dino_sprite[1][55][46] = 1;dino_sprite[1][55][47] = 1;dino_sprite[1][55][48] = 1;dino_sprite[1][55][49] = 1;dino_sprite[1][55][50] = 1;dino_sprite[1][55][51] = 1;dino_sprite[1][55][52] = 1;dino_sprite[1][55][53] = 1;dino_sprite[1][55][54] = 1;dino_sprite[1][55][55] = 1;dino_sprite[1][55][56] = 1;dino_sprite[1][55][57] = 1;dino_sprite[1][55][58] = 1;dino_sprite[1][55][59] = 1;dino_sprite[1][55][60] = 1;dino_sprite[1][55][61] = 1;dino_sprite[1][55][62] = 1;dino_sprite[1][55][63] = 1;dino_sprite[1][55][64] = 1;dino_sprite[1][55][65] = 1;dino_sprite[1][55][66] = 1;dino_sprite[1][55][67] = 1;dino_sprite[1][55][68] = 1;dino_sprite[1][55][69] = 1;dino_sprite[1][55][70] = 1;dino_sprite[1][55][71] = 1;dino_sprite[1][55][72] = 1;dino_sprite[1][55][73] = 1;dino_sprite[1][55][74] = 1;dino_sprite[1][55][75] = 1;dino_sprite[1][55][76] = 1;dino_sprite[1][55][77] = 1;dino_sprite[1][55][78] = 1;dino_sprite[1][55][79] = 1;dino_sprite[1][55][80] = 1;dino_sprite[1][55][81] = 1;dino_sprite[1][55][82] = 1;dino_sprite[1][55][83] = 1;dino_sprite[1][55][84] = 1;dino_sprite[1][55][85] = 1;dino_sprite[1][55][86] = 1;dino_sprite[1][55][87] = 1;dino_sprite[1][55][88] = 1;dino_sprite[1][55][89] = 1;dino_sprite[1][55][90] = 1;dino_sprite[1][55][91] = 1;dino_sprite[1][55][92] = 1;dino_sprite[1][55][93] = 1;dino_sprite[1][55][94] = 1;dino_sprite[1][55][95] = 1;dino_sprite[1][55][96] = 1;dino_sprite[1][55][97] = 1;dino_sprite[1][55][98] = 1;dino_sprite[1][55][99] = 1;dino_sprite[1][56][0] = 1;dino_sprite[1][56][1] = 1;dino_sprite[1][56][2] = 1;dino_sprite[1][56][3] = 1;dino_sprite[1][56][4] = 1;dino_sprite[1][56][5] = 1;dino_sprite[1][56][6] = 1;dino_sprite[1][56][7] = 1;dino_sprite[1][56][8] = 1;dino_sprite[1][56][9] = 1;dino_sprite[1][56][10] = 1;dino_sprite[1][56][11] = 1;dino_sprite[1][56][12] = 1;dino_sprite[1][56][13] = 1;dino_sprite[1][56][14] = 1;dino_sprite[1][56][15] = 1;dino_sprite[1][56][16] = 1;dino_sprite[1][56][17] = 1;dino_sprite[1][56][18] = 1;dino_sprite[1][56][19] = 1;dino_sprite[1][56][20] = 1;dino_sprite[1][56][21] = 1;dino_sprite[1][56][22] = 1;dino_sprite[1][56][23] = 1;dino_sprite[1][56][24] = 1;dino_sprite[1][56][25] = 1;dino_sprite[1][56][26] = 1;dino_sprite[1][56][27] = 1;dino_sprite[1][56][28] = 1;dino_sprite[1][56][29] = 1;dino_sprite[1][56][30] = 1;dino_sprite[1][56][31] = 1;dino_sprite[1][56][32] = 1;dino_sprite[1][56][33] = 1;dino_sprite[1][56][34] = 1;dino_sprite[1][56][35] = 1;dino_sprite[1][56][36] = 1;dino_sprite[1][56][37] = 1;dino_sprite[1][56][38] = 1;dino_sprite[1][56][39] = 1;dino_sprite[1][56][40] = 1;dino_sprite[1][56][41] = 1;dino_sprite[1][56][42] = 1;dino_sprite[1][56][43] = 1;dino_sprite[1][56][44] = 1;dino_sprite[1][56][45] = 1;dino_sprite[1][56][46] = 1;dino_sprite[1][56][47] = 1;dino_sprite[1][56][48] = 1;dino_sprite[1][56][49] = 1;dino_sprite[1][56][50] = 1;dino_sprite[1][56][51] = 1;dino_sprite[1][56][52] = 1;dino_sprite[1][56][53] = 1;dino_sprite[1][56][54] = 1;dino_sprite[1][56][55] = 1;dino_sprite[1][56][56] = 1;dino_sprite[1][56][57] = 1;dino_sprite[1][56][58] = 1;dino_sprite[1][56][59] = 1;dino_sprite[1][56][60] = 1;dino_sprite[1][56][61] = 1;dino_sprite[1][56][62] = 1;dino_sprite[1][56][63] = 1;dino_sprite[1][56][64] = 1;dino_sprite[1][56][65] = 1;dino_sprite[1][56][66] = 1;dino_sprite[1][56][67] = 1;dino_sprite[1][56][68] = 1;dino_sprite[1][56][69] = 1;dino_sprite[1][56][70] = 1;dino_sprite[1][56][71] = 1;dino_sprite[1][56][72] = 1;dino_sprite[1][56][73] = 1;dino_sprite[1][56][74] = 1;dino_sprite[1][56][75] = 1;dino_sprite[1][56][76] = 1;dino_sprite[1][56][77] = 1;dino_sprite[1][56][95] = 1;dino_sprite[1][56][96] = 1;dino_sprite[1][56][97] = 1;dino_sprite[1][56][98] = 1;dino_sprite[1][56][99] = 1;dino_sprite[1][57][0] = 1;dino_sprite[1][57][1] = 1;dino_sprite[1][57][2] = 1;dino_sprite[1][57][3] = 1;dino_sprite[1][57][4] = 1;dino_sprite[1][57][5] = 1;dino_sprite[1][57][6] = 1;dino_sprite[1][57][7] = 1;dino_sprite[1][57][8] = 1;dino_sprite[1][57][9] = 1;dino_sprite[1][57][10] = 1;dino_sprite[1][57][11] = 1;dino_sprite[1][57][12] = 1;dino_sprite[1][57][13] = 1;dino_sprite[1][57][14] = 1;dino_sprite[1][57][15] = 1;dino_sprite[1][57][16] = 1;dino_sprite[1][57][17] = 1;dino_sprite[1][57][18] = 1;dino_sprite[1][57][19] = 1;dino_sprite[1][57][20] = 1;dino_sprite[1][57][21] = 1;dino_sprite[1][57][22] = 1;dino_sprite[1][57][23] = 1;dino_sprite[1][57][24] = 1;dino_sprite[1][57][25] = 1;dino_sprite[1][57][26] = 1;dino_sprite[1][57][27] = 1;dino_sprite[1][57][28] = 1;dino_sprite[1][57][29] = 1;dino_sprite[1][57][30] = 1;dino_sprite[1][57][31] = 1;dino_sprite[1][57][32] = 1;dino_sprite[1][57][33] = 1;dino_sprite[1][57][34] = 1;dino_sprite[1][57][35] = 1;dino_sprite[1][57][36] = 1;dino_sprite[1][57][37] = 1;dino_sprite[1][57][38] = 1;dino_sprite[1][57][39] = 1;dino_sprite[1][57][40] = 1;dino_sprite[1][57][41] = 1;dino_sprite[1][57][42] = 1;dino_sprite[1][57][43] = 1;dino_sprite[1][57][44] = 1;dino_sprite[1][57][45] = 1;dino_sprite[1][57][46] = 1;dino_sprite[1][57][47] = 1;dino_sprite[1][57][48] = 1;dino_sprite[1][57][49] = 1;dino_sprite[1][57][50] = 1;dino_sprite[1][57][51] = 1;dino_sprite[1][57][52] = 1;dino_sprite[1][57][53] = 1;dino_sprite[1][57][54] = 1;dino_sprite[1][57][55] = 1;dino_sprite[1][57][56] = 1;dino_sprite[1][57][57] = 1;dino_sprite[1][57][58] = 1;dino_sprite[1][57][59] = 1;dino_sprite[1][57][60] = 1;dino_sprite[1][57][61] = 1;dino_sprite[1][57][62] = 1;dino_sprite[1][57][63] = 1;dino_sprite[1][57][64] = 1;dino_sprite[1][57][65] = 1;dino_sprite[1][57][66] = 1;dino_sprite[1][57][67] = 1;dino_sprite[1][57][68] = 1;dino_sprite[1][57][69] = 1;dino_sprite[1][57][70] = 1;dino_sprite[1][57][71] = 1;dino_sprite[1][57][72] = 1;dino_sprite[1][57][73] = 1;dino_sprite[1][57][74] = 1;dino_sprite[1][57][75] = 1;dino_sprite[1][57][76] = 1;dino_sprite[1][57][77] = 1;dino_sprite[1][57][95] = 1;dino_sprite[1][57][96] = 1;dino_sprite[1][57][97] = 1;dino_sprite[1][57][98] = 1;dino_sprite[1][57][99] = 1;dino_sprite[1][58][0] = 1;dino_sprite[1][58][1] = 1;dino_sprite[1][58][2] = 1;dino_sprite[1][58][3] = 1;dino_sprite[1][58][4] = 1;dino_sprite[1][58][5] = 1;dino_sprite[1][58][6] = 1;dino_sprite[1][58][7] = 1;dino_sprite[1][58][8] = 1;dino_sprite[1][58][9] = 1;dino_sprite[1][58][10] = 1;dino_sprite[1][58][11] = 1;dino_sprite[1][58][12] = 1;dino_sprite[1][58][13] = 1;dino_sprite[1][58][14] = 1;dino_sprite[1][58][15] = 1;dino_sprite[1][58][16] = 1;dino_sprite[1][58][17] = 1;dino_sprite[1][58][18] = 1;dino_sprite[1][58][19] = 1;dino_sprite[1][58][20] = 1;dino_sprite[1][58][21] = 1;dino_sprite[1][58][22] = 1;dino_sprite[1][58][23] = 1;dino_sprite[1][58][24] = 1;dino_sprite[1][58][25] = 1;dino_sprite[1][58][26] = 1;dino_sprite[1][58][27] = 1;dino_sprite[1][58][28] = 1;dino_sprite[1][58][29] = 1;dino_sprite[1][58][30] = 1;dino_sprite[1][58][31] = 1;dino_sprite[1][58][32] = 1;dino_sprite[1][58][33] = 1;dino_sprite[1][58][34] = 1;dino_sprite[1][58][35] = 1;dino_sprite[1][58][36] = 1;dino_sprite[1][58][37] = 1;dino_sprite[1][58][38] = 1;dino_sprite[1][58][39] = 1;dino_sprite[1][58][40] = 1;dino_sprite[1][58][41] = 1;dino_sprite[1][58][42] = 1;dino_sprite[1][58][43] = 1;dino_sprite[1][58][44] = 1;dino_sprite[1][58][45] = 1;dino_sprite[1][58][46] = 1;dino_sprite[1][58][47] = 1;dino_sprite[1][58][48] = 1;dino_sprite[1][58][49] = 1;dino_sprite[1][58][50] = 1;dino_sprite[1][58][51] = 1;dino_sprite[1][58][52] = 1;dino_sprite[1][58][53] = 1;dino_sprite[1][58][54] = 1;dino_sprite[1][58][55] = 1;dino_sprite[1][58][56] = 1;dino_sprite[1][58][57] = 1;dino_sprite[1][58][58] = 1;dino_sprite[1][58][59] = 1;dino_sprite[1][58][60] = 1;dino_sprite[1][58][61] = 1;dino_sprite[1][58][62] = 1;dino_sprite[1][58][63] = 1;dino_sprite[1][58][64] = 1;dino_sprite[1][58][65] = 1;dino_sprite[1][58][66] = 1;dino_sprite[1][58][67] = 1;dino_sprite[1][58][68] = 1;dino_sprite[1][58][69] = 1;dino_sprite[1][58][70] = 1;dino_sprite[1][58][71] = 1;dino_sprite[1][58][72] = 1;dino_sprite[1][58][73] = 1;dino_sprite[1][58][74] = 1;dino_sprite[1][58][75] = 1;dino_sprite[1][58][76] = 1;dino_sprite[1][58][77] = 1;dino_sprite[1][58][95] = 1;dino_sprite[1][58][96] = 1;dino_sprite[1][58][97] = 1;dino_sprite[1][58][98] = 1;dino_sprite[1][58][99] = 1;dino_sprite[1][59][0] = 1;dino_sprite[1][59][1] = 1;dino_sprite[1][59][2] = 1;dino_sprite[1][59][3] = 1;dino_sprite[1][59][4] = 1;dino_sprite[1][59][5] = 1;dino_sprite[1][59][6] = 1;dino_sprite[1][59][7] = 1;dino_sprite[1][59][8] = 1;dino_sprite[1][59][9] = 1;dino_sprite[1][59][10] = 1;dino_sprite[1][59][11] = 1;dino_sprite[1][59][12] = 1;dino_sprite[1][59][13] = 1;dino_sprite[1][59][14] = 1;dino_sprite[1][59][15] = 1;dino_sprite[1][59][16] = 1;dino_sprite[1][59][17] = 1;dino_sprite[1][59][18] = 1;dino_sprite[1][59][19] = 1;dino_sprite[1][59][20] = 1;dino_sprite[1][59][21] = 1;dino_sprite[1][59][22] = 1;dino_sprite[1][59][23] = 1;dino_sprite[1][59][24] = 1;dino_sprite[1][59][25] = 1;dino_sprite[1][59][26] = 1;dino_sprite[1][59][27] = 1;dino_sprite[1][59][28] = 1;dino_sprite[1][59][29] = 1;dino_sprite[1][59][30] = 1;dino_sprite[1][59][31] = 1;dino_sprite[1][59][32] = 1;dino_sprite[1][59][33] = 1;dino_sprite[1][59][34] = 1;dino_sprite[1][59][35] = 1;dino_sprite[1][59][36] = 1;dino_sprite[1][59][37] = 1;dino_sprite[1][59][38] = 1;dino_sprite[1][59][39] = 1;dino_sprite[1][59][40] = 1;dino_sprite[1][59][41] = 1;dino_sprite[1][59][42] = 1;dino_sprite[1][59][43] = 1;dino_sprite[1][59][44] = 1;dino_sprite[1][59][45] = 1;dino_sprite[1][59][46] = 1;dino_sprite[1][59][47] = 1;dino_sprite[1][59][48] = 1;dino_sprite[1][59][49] = 1;dino_sprite[1][59][50] = 1;dino_sprite[1][59][51] = 1;dino_sprite[1][59][52] = 1;dino_sprite[1][59][53] = 1;dino_sprite[1][59][54] = 1;dino_sprite[1][59][55] = 1;dino_sprite[1][59][56] = 1;dino_sprite[1][59][57] = 1;dino_sprite[1][59][58] = 1;dino_sprite[1][59][59] = 1;dino_sprite[1][59][60] = 1;dino_sprite[1][59][61] = 1;dino_sprite[1][59][62] = 1;dino_sprite[1][59][63] = 1;dino_sprite[1][59][64] = 1;dino_sprite[1][59][65] = 1;dino_sprite[1][59][66] = 1;dino_sprite[1][59][67] = 1;dino_sprite[1][59][68] = 1;dino_sprite[1][59][69] = 1;dino_sprite[1][59][70] = 1;dino_sprite[1][59][71] = 1;dino_sprite[1][59][72] = 1;dino_sprite[1][59][73] = 1;dino_sprite[1][59][74] = 1;dino_sprite[1][59][75] = 1;dino_sprite[1][59][76] = 1;dino_sprite[1][59][77] = 1;dino_sprite[1][59][95] = 1;dino_sprite[1][59][96] = 1;dino_sprite[1][59][97] = 1;dino_sprite[1][59][98] = 1;dino_sprite[1][59][99] = 1;dino_sprite[1][60][0] = 1;dino_sprite[1][60][1] = 1;dino_sprite[1][60][2] = 1;dino_sprite[1][60][3] = 1;dino_sprite[1][60][4] = 1;dino_sprite[1][60][5] = 1;dino_sprite[1][60][6] = 1;dino_sprite[1][60][7] = 1;dino_sprite[1][60][8] = 1;dino_sprite[1][60][9] = 1;dino_sprite[1][60][10] = 1;dino_sprite[1][60][11] = 1;dino_sprite[1][60][12] = 1;dino_sprite[1][60][13] = 1;dino_sprite[1][60][14] = 1;dino_sprite[1][60][15] = 1;dino_sprite[1][60][16] = 1;dino_sprite[1][60][17] = 1;dino_sprite[1][60][18] = 1;dino_sprite[1][60][19] = 1;dino_sprite[1][60][20] = 1;dino_sprite[1][60][21] = 1;dino_sprite[1][60][22] = 1;dino_sprite[1][60][23] = 1;dino_sprite[1][60][24] = 1;dino_sprite[1][60][25] = 1;dino_sprite[1][60][26] = 1;dino_sprite[1][60][27] = 1;dino_sprite[1][60][28] = 1;dino_sprite[1][60][29] = 1;dino_sprite[1][60][30] = 1;dino_sprite[1][60][31] = 1;dino_sprite[1][60][32] = 1;dino_sprite[1][60][33] = 1;dino_sprite[1][60][34] = 1;dino_sprite[1][60][35] = 1;dino_sprite[1][60][36] = 1;dino_sprite[1][60][37] = 1;dino_sprite[1][60][38] = 1;dino_sprite[1][60][39] = 1;dino_sprite[1][60][40] = 1;dino_sprite[1][60][41] = 1;dino_sprite[1][60][42] = 1;dino_sprite[1][60][43] = 1;dino_sprite[1][60][44] = 1;dino_sprite[1][60][45] = 1;dino_sprite[1][60][46] = 1;dino_sprite[1][60][47] = 1;dino_sprite[1][60][48] = 1;dino_sprite[1][60][49] = 1;dino_sprite[1][60][50] = 1;dino_sprite[1][60][51] = 1;dino_sprite[1][60][52] = 1;dino_sprite[1][60][53] = 1;dino_sprite[1][60][54] = 1;dino_sprite[1][60][55] = 1;dino_sprite[1][60][56] = 1;dino_sprite[1][60][57] = 1;dino_sprite[1][60][58] = 1;dino_sprite[1][60][59] = 1;dino_sprite[1][60][60] = 1;dino_sprite[1][60][61] = 1;dino_sprite[1][60][62] = 1;dino_sprite[1][60][63] = 1;dino_sprite[1][60][64] = 1;dino_sprite[1][60][65] = 1;dino_sprite[1][60][66] = 1;dino_sprite[1][60][67] = 1;dino_sprite[1][60][68] = 1;dino_sprite[1][60][69] = 1;dino_sprite[1][60][70] = 1;dino_sprite[1][60][71] = 1;dino_sprite[1][60][72] = 1;dino_sprite[1][60][73] = 1;dino_sprite[1][60][74] = 1;dino_sprite[1][60][75] = 1;dino_sprite[1][60][76] = 1;dino_sprite[1][60][77] = 1;dino_sprite[1][60][96] = 1;dino_sprite[1][60][97] = 1;dino_sprite[1][60][98] = 1;dino_sprite[1][60][99] = 1;dino_sprite[1][61][0] = 1;dino_sprite[1][61][1] = 1;dino_sprite[1][61][2] = 1;dino_sprite[1][61][3] = 1;dino_sprite[1][61][4] = 1;dino_sprite[1][61][5] = 1;dino_sprite[1][61][6] = 1;dino_sprite[1][61][10] = 1;dino_sprite[1][61][11] = 1;dino_sprite[1][61][12] = 1;dino_sprite[1][61][13] = 1;dino_sprite[1][61][14] = 1;dino_sprite[1][61][15] = 1;dino_sprite[1][61][16] = 1;dino_sprite[1][61][17] = 1;dino_sprite[1][61][18] = 1;dino_sprite[1][61][19] = 1;dino_sprite[1][61][20] = 1;dino_sprite[1][61][21] = 1;dino_sprite[1][61][22] = 1;dino_sprite[1][61][23] = 1;dino_sprite[1][61][24] = 1;dino_sprite[1][61][25] = 1;dino_sprite[1][61][26] = 1;dino_sprite[1][61][27] = 1;dino_sprite[1][61][28] = 1;dino_sprite[1][61][29] = 1;dino_sprite[1][61][30] = 1;dino_sprite[1][61][31] = 1;dino_sprite[1][61][32] = 1;dino_sprite[1][61][33] = 1;dino_sprite[1][61][34] = 1;dino_sprite[1][61][35] = 1;dino_sprite[1][61][36] = 1;dino_sprite[1][61][37] = 1;dino_sprite[1][61][38] = 1;dino_sprite[1][61][39] = 1;dino_sprite[1][61][40] = 1;dino_sprite[1][61][41] = 1;dino_sprite[1][61][42] = 1;dino_sprite[1][61][43] = 1;dino_sprite[1][61][44] = 1;dino_sprite[1][61][45] = 1;dino_sprite[1][61][46] = 1;dino_sprite[1][61][47] = 1;dino_sprite[1][61][48] = 1;dino_sprite[1][61][49] = 1;dino_sprite[1][61][50] = 1;dino_sprite[1][61][51] = 1;dino_sprite[1][61][52] = 1;dino_sprite[1][61][53] = 1;dino_sprite[1][61][54] = 1;dino_sprite[1][61][55] = 1;dino_sprite[1][61][56] = 1;dino_sprite[1][61][57] = 1;dino_sprite[1][61][58] = 1;dino_sprite[1][61][59] = 1;dino_sprite[1][61][60] = 1;dino_sprite[1][61][61] = 1;dino_sprite[1][61][62] = 1;dino_sprite[1][61][63] = 1;dino_sprite[1][61][64] = 1;dino_sprite[1][61][65] = 1;dino_sprite[1][61][66] = 1;dino_sprite[1][61][67] = 1;dino_sprite[1][61][68] = 1;dino_sprite[1][61][69] = 1;dino_sprite[1][61][70] = 1;dino_sprite[1][61][71] = 1;dino_sprite[1][61][72] = 1;dino_sprite[1][62][0] = 1;dino_sprite[1][62][1] = 1;dino_sprite[1][62][2] = 1;dino_sprite[1][62][3] = 1;dino_sprite[1][62][4] = 1;dino_sprite[1][62][5] = 1;dino_sprite[1][62][6] = 1;dino_sprite[1][62][10] = 1;dino_sprite[1][62][11] = 1;dino_sprite[1][62][12] = 1;dino_sprite[1][62][13] = 1;dino_sprite[1][62][14] = 1;dino_sprite[1][62][15] = 1;dino_sprite[1][62][16] = 1;dino_sprite[1][62][17] = 1;dino_sprite[1][62][18] = 1;dino_sprite[1][62][19] = 1;dino_sprite[1][62][20] = 1;dino_sprite[1][62][21] = 1;dino_sprite[1][62][22] = 1;dino_sprite[1][62][23] = 1;dino_sprite[1][62][24] = 1;dino_sprite[1][62][25] = 1;dino_sprite[1][62][26] = 1;dino_sprite[1][62][27] = 1;dino_sprite[1][62][28] = 1;dino_sprite[1][62][29] = 1;dino_sprite[1][62][30] = 1;dino_sprite[1][62][31] = 1;dino_sprite[1][62][32] = 1;dino_sprite[1][62][33] = 1;dino_sprite[1][62][34] = 1;dino_sprite[1][62][35] = 1;dino_sprite[1][62][36] = 1;dino_sprite[1][62][37] = 1;dino_sprite[1][62][38] = 1;dino_sprite[1][62][39] = 1;dino_sprite[1][62][40] = 1;dino_sprite[1][62][41] = 1;dino_sprite[1][62][42] = 1;dino_sprite[1][62][43] = 1;dino_sprite[1][62][44] = 1;dino_sprite[1][62][45] = 1;dino_sprite[1][62][46] = 1;dino_sprite[1][62][47] = 1;dino_sprite[1][62][48] = 1;dino_sprite[1][62][49] = 1;dino_sprite[1][62][50] = 1;dino_sprite[1][62][51] = 1;dino_sprite[1][62][52] = 1;dino_sprite[1][62][53] = 1;dino_sprite[1][62][54] = 1;dino_sprite[1][62][55] = 1;dino_sprite[1][62][56] = 1;dino_sprite[1][62][57] = 1;dino_sprite[1][62][58] = 1;dino_sprite[1][62][59] = 1;dino_sprite[1][62][60] = 1;dino_sprite[1][62][61] = 1;dino_sprite[1][62][62] = 1;dino_sprite[1][62][63] = 1;dino_sprite[1][62][64] = 1;dino_sprite[1][62][65] = 1;dino_sprite[1][62][66] = 1;dino_sprite[1][62][67] = 1;dino_sprite[1][62][68] = 1;dino_sprite[1][62][69] = 1;dino_sprite[1][62][70] = 1;dino_sprite[1][62][71] = 1;dino_sprite[1][62][72] = 1;dino_sprite[1][63][0] = 1;dino_sprite[1][63][1] = 1;dino_sprite[1][63][2] = 1;dino_sprite[1][63][3] = 1;dino_sprite[1][63][4] = 1;dino_sprite[1][63][5] = 1;dino_sprite[1][63][6] = 1;dino_sprite[1][63][10] = 1;dino_sprite[1][63][11] = 1;dino_sprite[1][63][12] = 1;dino_sprite[1][63][13] = 1;dino_sprite[1][63][14] = 1;dino_sprite[1][63][15] = 1;dino_sprite[1][63][16] = 1;dino_sprite[1][63][17] = 1;dino_sprite[1][63][18] = 1;dino_sprite[1][63][19] = 1;dino_sprite[1][63][20] = 1;dino_sprite[1][63][21] = 1;dino_sprite[1][63][22] = 1;dino_sprite[1][63][23] = 1;dino_sprite[1][63][24] = 1;dino_sprite[1][63][25] = 1;dino_sprite[1][63][26] = 1;dino_sprite[1][63][27] = 1;dino_sprite[1][63][28] = 1;dino_sprite[1][63][29] = 1;dino_sprite[1][63][30] = 1;dino_sprite[1][63][31] = 1;dino_sprite[1][63][32] = 1;dino_sprite[1][63][33] = 1;dino_sprite[1][63][34] = 1;dino_sprite[1][63][35] = 1;dino_sprite[1][63][36] = 1;dino_sprite[1][63][37] = 1;dino_sprite[1][63][38] = 1;dino_sprite[1][63][39] = 1;dino_sprite[1][63][40] = 1;dino_sprite[1][63][41] = 1;dino_sprite[1][63][42] = 1;dino_sprite[1][63][43] = 1;dino_sprite[1][63][44] = 1;dino_sprite[1][63][45] = 1;dino_sprite[1][63][46] = 1;dino_sprite[1][63][47] = 1;dino_sprite[1][63][48] = 1;dino_sprite[1][63][49] = 1;dino_sprite[1][63][50] = 1;dino_sprite[1][63][51] = 1;dino_sprite[1][63][52] = 1;dino_sprite[1][63][53] = 1;dino_sprite[1][63][54] = 1;dino_sprite[1][63][55] = 1;dino_sprite[1][63][56] = 1;dino_sprite[1][63][57] = 1;dino_sprite[1][63][58] = 1;dino_sprite[1][63][59] = 1;dino_sprite[1][63][60] = 1;dino_sprite[1][63][61] = 1;dino_sprite[1][63][62] = 1;dino_sprite[1][63][63] = 1;dino_sprite[1][63][64] = 1;dino_sprite[1][63][65] = 1;dino_sprite[1][63][66] = 1;dino_sprite[1][63][67] = 1;dino_sprite[1][63][68] = 1;dino_sprite[1][63][69] = 1;dino_sprite[1][63][70] = 1;dino_sprite[1][63][71] = 1;dino_sprite[1][63][72] = 1;dino_sprite[1][64][0] = 1;dino_sprite[1][64][1] = 1;dino_sprite[1][64][2] = 1;dino_sprite[1][64][3] = 1;dino_sprite[1][64][4] = 1;dino_sprite[1][64][5] = 1;dino_sprite[1][64][6] = 1;dino_sprite[1][64][10] = 1;dino_sprite[1][64][11] = 1;dino_sprite[1][64][12] = 1;dino_sprite[1][64][13] = 1;dino_sprite[1][64][14] = 1;dino_sprite[1][64][15] = 1;dino_sprite[1][64][16] = 1;dino_sprite[1][64][17] = 1;dino_sprite[1][64][18] = 1;dino_sprite[1][64][19] = 1;dino_sprite[1][64][20] = 1;dino_sprite[1][64][21] = 1;dino_sprite[1][64][22] = 1;dino_sprite[1][64][23] = 1;dino_sprite[1][64][24] = 1;dino_sprite[1][64][25] = 1;dino_sprite[1][64][26] = 1;dino_sprite[1][64][27] = 1;dino_sprite[1][64][28] = 1;dino_sprite[1][64][29] = 1;dino_sprite[1][64][30] = 1;dino_sprite[1][64][31] = 1;dino_sprite[1][64][32] = 1;dino_sprite[1][64][33] = 1;dino_sprite[1][64][34] = 1;dino_sprite[1][64][35] = 1;dino_sprite[1][64][36] = 1;dino_sprite[1][64][37] = 1;dino_sprite[1][64][38] = 1;dino_sprite[1][64][39] = 1;dino_sprite[1][64][40] = 1;dino_sprite[1][64][41] = 1;dino_sprite[1][64][42] = 1;dino_sprite[1][64][43] = 1;dino_sprite[1][64][44] = 1;dino_sprite[1][64][45] = 1;dino_sprite[1][64][46] = 1;dino_sprite[1][64][47] = 1;dino_sprite[1][64][48] = 1;dino_sprite[1][64][49] = 1;dino_sprite[1][64][50] = 1;dino_sprite[1][64][51] = 1;dino_sprite[1][64][52] = 1;dino_sprite[1][64][53] = 1;dino_sprite[1][64][54] = 1;dino_sprite[1][64][55] = 1;dino_sprite[1][64][56] = 1;dino_sprite[1][64][57] = 1;dino_sprite[1][64][58] = 1;dino_sprite[1][64][59] = 1;dino_sprite[1][64][60] = 1;dino_sprite[1][64][61] = 1;dino_sprite[1][64][62] = 1;dino_sprite[1][64][63] = 1;dino_sprite[1][64][64] = 1;dino_sprite[1][64][65] = 1;dino_sprite[1][64][66] = 1;dino_sprite[1][64][67] = 1;dino_sprite[1][64][68] = 1;dino_sprite[1][64][69] = 1;dino_sprite[1][64][70] = 1;dino_sprite[1][64][71] = 1;dino_sprite[1][64][72] = 1;dino_sprite[1][65][0] = 1;dino_sprite[1][65][1] = 1;dino_sprite[1][65][2] = 1;dino_sprite[1][65][3] = 1;dino_sprite[1][65][4] = 1;dino_sprite[1][65][5] = 1;dino_sprite[1][65][6] = 1;dino_sprite[1][65][8] = 1;dino_sprite[1][65][10] = 1;dino_sprite[1][65][11] = 1;dino_sprite[1][65][12] = 1;dino_sprite[1][65][13] = 1;dino_sprite[1][65][14] = 1;dino_sprite[1][65][15] = 1;dino_sprite[1][65][16] = 1;dino_sprite[1][65][17] = 1;dino_sprite[1][65][18] = 1;dino_sprite[1][65][19] = 1;dino_sprite[1][65][20] = 1;dino_sprite[1][65][21] = 1;dino_sprite[1][65][22] = 1;dino_sprite[1][65][23] = 1;dino_sprite[1][65][24] = 1;dino_sprite[1][65][25] = 1;dino_sprite[1][65][26] = 1;dino_sprite[1][65][27] = 1;dino_sprite[1][65][28] = 1;dino_sprite[1][65][29] = 1;dino_sprite[1][65][30] = 1;dino_sprite[1][65][31] = 1;dino_sprite[1][65][32] = 1;dino_sprite[1][65][33] = 1;dino_sprite[1][65][34] = 1;dino_sprite[1][65][35] = 1;dino_sprite[1][65][36] = 1;dino_sprite[1][65][37] = 1;dino_sprite[1][65][38] = 1;dino_sprite[1][65][39] = 1;dino_sprite[1][65][40] = 1;dino_sprite[1][65][41] = 1;dino_sprite[1][65][42] = 1;dino_sprite[1][65][43] = 1;dino_sprite[1][65][44] = 1;dino_sprite[1][65][45] = 1;dino_sprite[1][65][46] = 1;dino_sprite[1][65][47] = 1;dino_sprite[1][65][48] = 1;dino_sprite[1][65][49] = 1;dino_sprite[1][65][50] = 1;dino_sprite[1][65][51] = 1;dino_sprite[1][65][52] = 1;dino_sprite[1][65][53] = 1;dino_sprite[1][65][54] = 1;dino_sprite[1][65][55] = 1;dino_sprite[1][65][56] = 1;dino_sprite[1][65][57] = 1;dino_sprite[1][65][58] = 1;dino_sprite[1][65][59] = 1;dino_sprite[1][65][60] = 1;dino_sprite[1][65][61] = 1;dino_sprite[1][65][62] = 1;dino_sprite[1][65][63] = 1;dino_sprite[1][65][64] = 1;dino_sprite[1][65][65] = 1;dino_sprite[1][65][66] = 1;dino_sprite[1][65][67] = 1;dino_sprite[1][65][68] = 1;dino_sprite[1][65][69] = 1;dino_sprite[1][65][70] = 1;dino_sprite[1][65][71] = 1;dino_sprite[1][65][72] = 1;dino_sprite[1][66][0] = 1;dino_sprite[1][66][1] = 1;dino_sprite[1][66][2] = 1;dino_sprite[1][66][3] = 1;dino_sprite[1][66][4] = 1;dino_sprite[1][66][5] = 1;dino_sprite[1][66][6] = 1;dino_sprite[1][66][7] = 1;dino_sprite[1][66][8] = 1;dino_sprite[1][66][9] = 1;dino_sprite[1][66][10] = 1;dino_sprite[1][66][11] = 1;dino_sprite[1][66][12] = 1;dino_sprite[1][66][13] = 1;dino_sprite[1][66][14] = 1;dino_sprite[1][66][15] = 1;dino_sprite[1][66][16] = 1;dino_sprite[1][66][17] = 1;dino_sprite[1][66][18] = 1;dino_sprite[1][66][19] = 1;dino_sprite[1][66][20] = 1;dino_sprite[1][66][21] = 1;dino_sprite[1][66][22] = 1;dino_sprite[1][66][23] = 1;dino_sprite[1][66][24] = 1;dino_sprite[1][66][25] = 1;dino_sprite[1][66][26] = 1;dino_sprite[1][66][27] = 1;dino_sprite[1][66][28] = 1;dino_sprite[1][66][29] = 1;dino_sprite[1][66][30] = 1;dino_sprite[1][66][31] = 1;dino_sprite[1][66][32] = 1;dino_sprite[1][66][33] = 1;dino_sprite[1][66][34] = 1;dino_sprite[1][66][35] = 1;dino_sprite[1][66][36] = 1;dino_sprite[1][66][37] = 1;dino_sprite[1][66][38] = 1;dino_sprite[1][66][39] = 1;dino_sprite[1][66][40] = 1;dino_sprite[1][66][41] = 1;dino_sprite[1][66][42] = 1;dino_sprite[1][66][43] = 1;dino_sprite[1][66][44] = 1;dino_sprite[1][66][45] = 1;dino_sprite[1][66][46] = 1;dino_sprite[1][66][47] = 1;dino_sprite[1][66][48] = 1;dino_sprite[1][66][49] = 1;dino_sprite[1][66][50] = 1;dino_sprite[1][66][51] = 1;dino_sprite[1][66][52] = 1;dino_sprite[1][66][53] = 1;dino_sprite[1][66][54] = 1;dino_sprite[1][66][55] = 1;dino_sprite[1][66][56] = 1;dino_sprite[1][66][57] = 1;dino_sprite[1][66][58] = 1;dino_sprite[1][66][59] = 1;dino_sprite[1][66][60] = 1;dino_sprite[1][66][61] = 1;dino_sprite[1][66][62] = 1;dino_sprite[1][66][63] = 1;dino_sprite[1][66][64] = 1;dino_sprite[1][66][65] = 1;dino_sprite[1][67][0] = 1;dino_sprite[1][67][1] = 1;dino_sprite[1][67][2] = 1;dino_sprite[1][67][3] = 1;dino_sprite[1][67][4] = 1;dino_sprite[1][67][5] = 1;dino_sprite[1][67][6] = 1;dino_sprite[1][67][7] = 1;dino_sprite[1][67][8] = 1;dino_sprite[1][67][9] = 1;dino_sprite[1][67][10] = 1;dino_sprite[1][67][11] = 1;dino_sprite[1][67][12] = 1;dino_sprite[1][67][13] = 1;dino_sprite[1][67][14] = 1;dino_sprite[1][67][15] = 1;dino_sprite[1][67][16] = 1;dino_sprite[1][67][17] = 1;dino_sprite[1][67][18] = 1;dino_sprite[1][67][19] = 1;dino_sprite[1][67][20] = 1;dino_sprite[1][67][21] = 1;dino_sprite[1][67][22] = 1;dino_sprite[1][67][23] = 1;dino_sprite[1][67][24] = 1;dino_sprite[1][67][25] = 1;dino_sprite[1][67][26] = 1;dino_sprite[1][67][27] = 1;dino_sprite[1][67][28] = 1;dino_sprite[1][67][29] = 1;dino_sprite[1][67][30] = 1;dino_sprite[1][67][31] = 1;dino_sprite[1][67][32] = 1;dino_sprite[1][67][33] = 1;dino_sprite[1][67][34] = 1;dino_sprite[1][67][35] = 1;dino_sprite[1][67][36] = 1;dino_sprite[1][67][37] = 1;dino_sprite[1][67][38] = 1;dino_sprite[1][67][39] = 1;dino_sprite[1][67][40] = 1;dino_sprite[1][67][41] = 1;dino_sprite[1][67][42] = 1;dino_sprite[1][67][43] = 1;dino_sprite[1][67][44] = 1;dino_sprite[1][67][45] = 1;dino_sprite[1][67][46] = 1;dino_sprite[1][67][47] = 1;dino_sprite[1][67][48] = 1;dino_sprite[1][67][49] = 1;dino_sprite[1][67][50] = 1;dino_sprite[1][67][51] = 1;dino_sprite[1][67][52] = 1;dino_sprite[1][67][53] = 1;dino_sprite[1][67][54] = 1;dino_sprite[1][67][55] = 1;dino_sprite[1][67][56] = 1;dino_sprite[1][67][57] = 1;dino_sprite[1][67][58] = 1;dino_sprite[1][67][59] = 1;dino_sprite[1][67][60] = 1;dino_sprite[1][67][61] = 1;dino_sprite[1][67][62] = 1;dino_sprite[1][67][63] = 1;dino_sprite[1][67][64] = 1;dino_sprite[1][67][65] = 1;dino_sprite[1][68][0] = 1;dino_sprite[1][68][1] = 1;dino_sprite[1][68][2] = 1;dino_sprite[1][68][3] = 1;dino_sprite[1][68][4] = 1;dino_sprite[1][68][5] = 1;dino_sprite[1][68][6] = 1;dino_sprite[1][68][7] = 1;dino_sprite[1][68][8] = 1;dino_sprite[1][68][9] = 1;dino_sprite[1][68][10] = 1;dino_sprite[1][68][11] = 1;dino_sprite[1][68][12] = 1;dino_sprite[1][68][13] = 1;dino_sprite[1][68][14] = 1;dino_sprite[1][68][15] = 1;dino_sprite[1][68][16] = 1;dino_sprite[1][68][17] = 1;dino_sprite[1][68][18] = 1;dino_sprite[1][68][19] = 1;dino_sprite[1][68][20] = 1;dino_sprite[1][68][21] = 1;dino_sprite[1][68][22] = 1;dino_sprite[1][68][23] = 1;dino_sprite[1][68][24] = 1;dino_sprite[1][68][25] = 1;dino_sprite[1][68][26] = 1;dino_sprite[1][68][27] = 1;dino_sprite[1][68][28] = 1;dino_sprite[1][68][29] = 1;dino_sprite[1][68][30] = 1;dino_sprite[1][68][31] = 1;dino_sprite[1][68][32] = 1;dino_sprite[1][68][33] = 1;dino_sprite[1][68][34] = 1;dino_sprite[1][68][35] = 1;dino_sprite[1][68][36] = 1;dino_sprite[1][68][37] = 1;dino_sprite[1][68][38] = 1;dino_sprite[1][68][39] = 1;dino_sprite[1][68][40] = 1;dino_sprite[1][68][41] = 1;dino_sprite[1][68][42] = 1;dino_sprite[1][68][43] = 1;dino_sprite[1][68][44] = 1;dino_sprite[1][68][45] = 1;dino_sprite[1][68][46] = 1;dino_sprite[1][68][47] = 1;dino_sprite[1][68][48] = 1;dino_sprite[1][68][49] = 1;dino_sprite[1][68][50] = 1;dino_sprite[1][68][51] = 1;dino_sprite[1][68][52] = 1;dino_sprite[1][68][53] = 1;dino_sprite[1][68][54] = 1;dino_sprite[1][68][55] = 1;dino_sprite[1][68][56] = 1;dino_sprite[1][68][57] = 1;dino_sprite[1][68][58] = 1;dino_sprite[1][68][59] = 1;dino_sprite[1][68][60] = 1;dino_sprite[1][68][61] = 1;dino_sprite[1][68][62] = 1;dino_sprite[1][68][63] = 1;dino_sprite[1][68][64] = 1;dino_sprite[1][68][65] = 1;dino_sprite[1][69][0] = 1;dino_sprite[1][69][1] = 1;dino_sprite[1][69][2] = 1;dino_sprite[1][69][3] = 1;dino_sprite[1][69][4] = 1;dino_sprite[1][69][5] = 1;dino_sprite[1][69][6] = 1;dino_sprite[1][69][7] = 1;dino_sprite[1][69][8] = 1;dino_sprite[1][69][9] = 1;dino_sprite[1][69][10] = 1;dino_sprite[1][69][11] = 1;dino_sprite[1][69][12] = 1;dino_sprite[1][69][13] = 1;dino_sprite[1][69][14] = 1;dino_sprite[1][69][15] = 1;dino_sprite[1][69][16] = 1;dino_sprite[1][69][17] = 1;dino_sprite[1][69][18] = 1;dino_sprite[1][69][19] = 1;dino_sprite[1][69][20] = 1;dino_sprite[1][69][21] = 1;dino_sprite[1][69][22] = 1;dino_sprite[1][69][23] = 1;dino_sprite[1][69][24] = 1;dino_sprite[1][69][25] = 1;dino_sprite[1][69][26] = 1;dino_sprite[1][69][27] = 1;dino_sprite[1][69][28] = 1;dino_sprite[1][69][29] = 1;dino_sprite[1][69][30] = 1;dino_sprite[1][69][31] = 1;dino_sprite[1][69][32] = 1;dino_sprite[1][69][33] = 1;dino_sprite[1][69][34] = 1;dino_sprite[1][69][35] = 1;dino_sprite[1][69][36] = 1;dino_sprite[1][69][37] = 1;dino_sprite[1][69][38] = 1;dino_sprite[1][69][39] = 1;dino_sprite[1][69][40] = 1;dino_sprite[1][69][41] = 1;dino_sprite[1][69][42] = 1;dino_sprite[1][69][43] = 1;dino_sprite[1][69][44] = 1;dino_sprite[1][69][45] = 1;dino_sprite[1][69][46] = 1;dino_sprite[1][69][47] = 1;dino_sprite[1][69][48] = 1;dino_sprite[1][69][49] = 1;dino_sprite[1][69][50] = 1;dino_sprite[1][69][51] = 1;dino_sprite[1][69][52] = 1;dino_sprite[1][69][53] = 1;dino_sprite[1][69][54] = 1;dino_sprite[1][69][55] = 1;dino_sprite[1][69][56] = 1;dino_sprite[1][69][57] = 1;dino_sprite[1][69][58] = 1;dino_sprite[1][69][59] = 1;dino_sprite[1][69][60] = 1;dino_sprite[1][69][61] = 1;dino_sprite[1][69][62] = 1;dino_sprite[1][69][63] = 1;dino_sprite[1][69][64] = 1;dino_sprite[1][69][65] = 1;dino_sprite[1][70][0] = 1;dino_sprite[1][70][1] = 1;dino_sprite[1][70][2] = 1;dino_sprite[1][70][3] = 1;dino_sprite[1][70][4] = 1;dino_sprite[1][70][5] = 1;dino_sprite[1][70][6] = 1;dino_sprite[1][70][7] = 1;dino_sprite[1][70][8] = 1;dino_sprite[1][70][9] = 1;dino_sprite[1][70][10] = 1;dino_sprite[1][70][11] = 1;dino_sprite[1][70][12] = 1;dino_sprite[1][70][13] = 1;dino_sprite[1][70][14] = 1;dino_sprite[1][70][15] = 1;dino_sprite[1][70][16] = 1;dino_sprite[1][70][17] = 1;dino_sprite[1][70][18] = 1;dino_sprite[1][70][19] = 1;dino_sprite[1][70][20] = 1;dino_sprite[1][70][21] = 1;dino_sprite[1][70][22] = 1;dino_sprite[1][70][23] = 1;dino_sprite[1][70][24] = 1;dino_sprite[1][70][25] = 1;dino_sprite[1][70][26] = 1;dino_sprite[1][70][27] = 1;dino_sprite[1][70][28] = 1;dino_sprite[1][70][29] = 1;dino_sprite[1][70][30] = 1;dino_sprite[1][70][31] = 1;dino_sprite[1][70][32] = 1;dino_sprite[1][70][33] = 1;dino_sprite[1][70][34] = 1;dino_sprite[1][70][35] = 1;dino_sprite[1][70][36] = 1;dino_sprite[1][70][37] = 1;dino_sprite[1][70][38] = 1;dino_sprite[1][70][39] = 1;dino_sprite[1][70][40] = 1;dino_sprite[1][70][41] = 1;dino_sprite[1][70][42] = 1;dino_sprite[1][70][43] = 1;dino_sprite[1][70][44] = 1;dino_sprite[1][70][45] = 1;dino_sprite[1][70][46] = 1;dino_sprite[1][70][47] = 1;dino_sprite[1][70][48] = 1;dino_sprite[1][70][49] = 1;dino_sprite[1][70][50] = 1;dino_sprite[1][70][51] = 1;dino_sprite[1][70][52] = 1;dino_sprite[1][70][53] = 1;dino_sprite[1][70][54] = 1;dino_sprite[1][70][55] = 1;dino_sprite[1][70][56] = 1;dino_sprite[1][70][57] = 1;dino_sprite[1][70][58] = 1;dino_sprite[1][70][59] = 1;dino_sprite[1][70][60] = 1;dino_sprite[1][70][61] = 1;dino_sprite[1][70][62] = 1;dino_sprite[1][70][63] = 1;dino_sprite[1][70][64] = 1;dino_sprite[1][70][65] = 1;dino_sprite[1][71][0] = 1;dino_sprite[1][71][1] = 1;dino_sprite[1][71][2] = 1;dino_sprite[1][71][3] = 1;dino_sprite[1][71][4] = 1;dino_sprite[1][71][5] = 1;dino_sprite[1][71][6] = 1;dino_sprite[1][71][7] = 1;dino_sprite[1][71][8] = 1;dino_sprite[1][71][9] = 1;dino_sprite[1][71][10] = 1;dino_sprite[1][71][11] = 1;dino_sprite[1][71][12] = 1;dino_sprite[1][71][13] = 1;dino_sprite[1][71][14] = 1;dino_sprite[1][71][15] = 1;dino_sprite[1][71][16] = 1;dino_sprite[1][71][17] = 1;dino_sprite[1][71][18] = 1;dino_sprite[1][71][19] = 1;dino_sprite[1][71][20] = 1;dino_sprite[1][71][21] = 1;dino_sprite[1][71][22] = 1;dino_sprite[1][71][23] = 1;dino_sprite[1][71][24] = 1;dino_sprite[1][71][25] = 1;dino_sprite[1][71][26] = 1;dino_sprite[1][71][27] = 1;dino_sprite[1][71][28] = 1;dino_sprite[1][71][29] = 1;dino_sprite[1][71][30] = 1;dino_sprite[1][71][31] = 1;dino_sprite[1][71][32] = 1;dino_sprite[1][71][33] = 1;dino_sprite[1][71][34] = 1;dino_sprite[1][71][35] = 1;dino_sprite[1][71][36] = 1;dino_sprite[1][71][37] = 1;dino_sprite[1][71][38] = 1;dino_sprite[1][71][39] = 1;dino_sprite[1][71][40] = 1;dino_sprite[1][71][41] = 1;dino_sprite[1][71][43] = 1;dino_sprite[1][71][44] = 1;dino_sprite[1][71][45] = 1;dino_sprite[1][71][46] = 1;dino_sprite[1][71][47] = 1;dino_sprite[1][71][48] = 1;dino_sprite[1][71][49] = 1;dino_sprite[1][72][0] = 1;dino_sprite[1][72][1] = 1;dino_sprite[1][72][2] = 1;dino_sprite[1][72][3] = 1;dino_sprite[1][72][4] = 1;dino_sprite[1][72][5] = 1;dino_sprite[1][72][6] = 1;dino_sprite[1][72][7] = 1;dino_sprite[1][72][8] = 1;dino_sprite[1][72][9] = 1;dino_sprite[1][72][10] = 1;dino_sprite[1][72][11] = 1;dino_sprite[1][72][12] = 1;dino_sprite[1][72][13] = 1;dino_sprite[1][72][14] = 1;dino_sprite[1][72][15] = 1;dino_sprite[1][72][16] = 1;dino_sprite[1][72][17] = 1;dino_sprite[1][72][18] = 1;dino_sprite[1][72][19] = 1;dino_sprite[1][72][20] = 1;dino_sprite[1][72][21] = 1;dino_sprite[1][72][22] = 1;dino_sprite[1][72][23] = 1;dino_sprite[1][72][24] = 1;dino_sprite[1][72][25] = 1;dino_sprite[1][72][26] = 1;dino_sprite[1][72][27] = 1;dino_sprite[1][72][28] = 1;dino_sprite[1][72][29] = 1;dino_sprite[1][72][30] = 1;dino_sprite[1][72][31] = 1;dino_sprite[1][72][32] = 1;dino_sprite[1][72][33] = 1;dino_sprite[1][72][34] = 1;dino_sprite[1][72][35] = 1;dino_sprite[1][72][43] = 1;dino_sprite[1][72][44] = 1;dino_sprite[1][72][45] = 1;dino_sprite[1][72][46] = 1;dino_sprite[1][72][47] = 1;dino_sprite[1][72][48] = 1;dino_sprite[1][72][49] = 1;dino_sprite[1][73][0] = 1;dino_sprite[1][73][1] = 1;dino_sprite[1][73][2] = 1;dino_sprite[1][73][3] = 1;dino_sprite[1][73][4] = 1;dino_sprite[1][73][5] = 1;dino_sprite[1][73][6] = 1;dino_sprite[1][73][7] = 1;dino_sprite[1][73][8] = 1;dino_sprite[1][73][9] = 1;dino_sprite[1][73][10] = 1;dino_sprite[1][73][11] = 1;dino_sprite[1][73][12] = 1;dino_sprite[1][73][13] = 1;dino_sprite[1][73][14] = 1;dino_sprite[1][73][15] = 1;dino_sprite[1][73][16] = 1;dino_sprite[1][73][17] = 1;dino_sprite[1][73][18] = 1;dino_sprite[1][73][19] = 1;dino_sprite[1][73][20] = 1;dino_sprite[1][73][21] = 1;dino_sprite[1][73][22] = 1;dino_sprite[1][73][23] = 1;dino_sprite[1][73][24] = 1;dino_sprite[1][73][25] = 1;dino_sprite[1][73][26] = 1;dino_sprite[1][73][27] = 1;dino_sprite[1][73][28] = 1;dino_sprite[1][73][29] = 1;dino_sprite[1][73][30] = 1;dino_sprite[1][73][31] = 1;dino_sprite[1][73][32] = 1;dino_sprite[1][73][33] = 1;dino_sprite[1][73][34] = 1;dino_sprite[1][73][35] = 1;dino_sprite[1][73][43] = 1;dino_sprite[1][73][44] = 1;dino_sprite[1][73][45] = 1;dino_sprite[1][73][46] = 1;dino_sprite[1][73][47] = 1;dino_sprite[1][73][48] = 1;dino_sprite[1][73][49] = 1;dino_sprite[1][74][0] = 1;dino_sprite[1][74][1] = 1;dino_sprite[1][74][2] = 1;dino_sprite[1][74][3] = 1;dino_sprite[1][74][4] = 1;dino_sprite[1][74][5] = 1;dino_sprite[1][74][6] = 1;dino_sprite[1][74][7] = 1;dino_sprite[1][74][8] = 1;dino_sprite[1][74][9] = 1;dino_sprite[1][74][10] = 1;dino_sprite[1][74][11] = 1;dino_sprite[1][74][12] = 1;dino_sprite[1][74][13] = 1;dino_sprite[1][74][14] = 1;dino_sprite[1][74][15] = 1;dino_sprite[1][74][16] = 1;dino_sprite[1][74][17] = 1;dino_sprite[1][74][18] = 1;dino_sprite[1][74][19] = 1;dino_sprite[1][74][20] = 1;dino_sprite[1][74][21] = 1;dino_sprite[1][74][22] = 1;dino_sprite[1][74][23] = 1;dino_sprite[1][74][24] = 1;dino_sprite[1][74][25] = 1;dino_sprite[1][74][26] = 1;dino_sprite[1][74][27] = 1;dino_sprite[1][74][28] = 1;dino_sprite[1][74][29] = 1;dino_sprite[1][74][30] = 1;dino_sprite[1][74][31] = 1;dino_sprite[1][74][32] = 1;dino_sprite[1][74][33] = 1;dino_sprite[1][74][34] = 1;dino_sprite[1][74][35] = 1;dino_sprite[1][74][43] = 1;dino_sprite[1][74][44] = 1;dino_sprite[1][74][45] = 1;dino_sprite[1][74][46] = 1;dino_sprite[1][74][47] = 1;dino_sprite[1][74][48] = 1;dino_sprite[1][74][49] = 1;dino_sprite[1][75][0] = 1;dino_sprite[1][75][1] = 1;dino_sprite[1][75][2] = 1;dino_sprite[1][75][3] = 1;dino_sprite[1][75][4] = 1;dino_sprite[1][75][5] = 1;dino_sprite[1][75][6] = 1;dino_sprite[1][75][7] = 1;dino_sprite[1][75][8] = 1;dino_sprite[1][75][9] = 1;dino_sprite[1][75][10] = 1;dino_sprite[1][75][11] = 1;dino_sprite[1][75][12] = 1;dino_sprite[1][75][13] = 1;dino_sprite[1][75][14] = 1;dino_sprite[1][75][15] = 1;dino_sprite[1][75][16] = 1;dino_sprite[1][75][17] = 1;dino_sprite[1][75][18] = 1;dino_sprite[1][75][19] = 1;dino_sprite[1][75][20] = 1;dino_sprite[1][75][21] = 1;dino_sprite[1][75][22] = 1;dino_sprite[1][75][23] = 1;dino_sprite[1][75][24] = 1;dino_sprite[1][75][25] = 1;dino_sprite[1][75][26] = 1;dino_sprite[1][75][27] = 1;dino_sprite[1][75][28] = 1;dino_sprite[1][75][29] = 1;dino_sprite[1][75][30] = 1;dino_sprite[1][75][31] = 1;dino_sprite[1][75][32] = 1;dino_sprite[1][75][33] = 1;dino_sprite[1][75][34] = 1;dino_sprite[1][75][35] = 1;dino_sprite[1][75][43] = 1;dino_sprite[1][75][44] = 1;dino_sprite[1][75][45] = 1;dino_sprite[1][75][46] = 1;dino_sprite[1][75][47] = 1;dino_sprite[1][75][48] = 1;dino_sprite[1][75][49] = 1;dino_sprite[1][75][50] = 1;dino_sprite[1][75][51] = 1;dino_sprite[1][75][52] = 1;dino_sprite[1][75][53] = 1;dino_sprite[1][75][54] = 1;dino_sprite[1][76][0] = 1;dino_sprite[1][76][1] = 1;dino_sprite[1][76][2] = 1;dino_sprite[1][76][3] = 1;dino_sprite[1][76][4] = 1;dino_sprite[1][76][5] = 1;dino_sprite[1][76][6] = 1;dino_sprite[1][76][7] = 1;dino_sprite[1][76][8] = 1;dino_sprite[1][76][9] = 1;dino_sprite[1][76][10] = 1;dino_sprite[1][76][11] = 1;dino_sprite[1][76][12] = 1;dino_sprite[1][76][13] = 1;dino_sprite[1][76][14] = 1;dino_sprite[1][76][15] = 1;dino_sprite[1][76][16] = 1;dino_sprite[1][76][17] = 1;dino_sprite[1][76][18] = 1;dino_sprite[1][76][19] = 1;dino_sprite[1][76][20] = 1;dino_sprite[1][76][21] = 1;dino_sprite[1][76][22] = 1;dino_sprite[1][76][23] = 1;dino_sprite[1][76][24] = 1;dino_sprite[1][76][25] = 1;dino_sprite[1][76][26] = 1;dino_sprite[1][76][27] = 1;dino_sprite[1][76][28] = 1;dino_sprite[1][76][29] = 1;dino_sprite[1][76][30] = 1;dino_sprite[1][76][31] = 1;dino_sprite[1][76][32] = 1;dino_sprite[1][76][33] = 1;dino_sprite[1][76][34] = 1;dino_sprite[1][76][35] = 1;dino_sprite[1][76][43] = 1;dino_sprite[1][76][44] = 1;dino_sprite[1][76][45] = 1;dino_sprite[1][76][46] = 1;dino_sprite[1][76][47] = 1;dino_sprite[1][76][48] = 1;dino_sprite[1][76][49] = 1;dino_sprite[1][76][50] = 1;dino_sprite[1][76][51] = 1;dino_sprite[1][76][52] = 1;dino_sprite[1][76][53] = 1;dino_sprite[1][76][54] = 1;dino_sprite[1][77][0] = 1;dino_sprite[1][77][1] = 1;dino_sprite[1][77][2] = 1;dino_sprite[1][77][3] = 1;dino_sprite[1][77][4] = 1;dino_sprite[1][77][5] = 1;dino_sprite[1][77][6] = 1;dino_sprite[1][77][7] = 1;dino_sprite[1][77][8] = 1;dino_sprite[1][77][9] = 1;dino_sprite[1][77][10] = 1;dino_sprite[1][77][11] = 1;dino_sprite[1][77][12] = 1;dino_sprite[1][77][13] = 1;dino_sprite[1][77][14] = 1;dino_sprite[1][77][15] = 1;dino_sprite[1][77][16] = 1;dino_sprite[1][77][17] = 1;dino_sprite[1][77][18] = 1;dino_sprite[1][77][19] = 1;dino_sprite[1][77][20] = 1;dino_sprite[1][77][21] = 1;dino_sprite[1][77][22] = 1;dino_sprite[1][77][23] = 1;dino_sprite[1][77][24] = 1;dino_sprite[1][77][25] = 1;dino_sprite[1][77][29] = 1;dino_sprite[1][77][30] = 1;dino_sprite[1][77][31] = 1;dino_sprite[1][77][32] = 1;dino_sprite[1][77][33] = 1;dino_sprite[1][77][34] = 1;dino_sprite[1][77][35] = 1;dino_sprite[1][77][43] = 1;dino_sprite[1][77][44] = 1;dino_sprite[1][77][45] = 1;dino_sprite[1][77][46] = 1;dino_sprite[1][77][47] = 1;dino_sprite[1][77][48] = 1;dino_sprite[1][77][49] = 1;dino_sprite[1][77][50] = 1;dino_sprite[1][77][51] = 1;dino_sprite[1][77][52] = 1;dino_sprite[1][77][53] = 1;dino_sprite[1][77][54] = 1;dino_sprite[1][78][0] = 1;dino_sprite[1][78][1] = 1;dino_sprite[1][78][2] = 1;dino_sprite[1][78][3] = 1;dino_sprite[1][78][4] = 1;dino_sprite[1][78][5] = 1;dino_sprite[1][78][6] = 1;dino_sprite[1][78][7] = 1;dino_sprite[1][78][8] = 1;dino_sprite[1][78][9] = 1;dino_sprite[1][78][10] = 1;dino_sprite[1][78][11] = 1;dino_sprite[1][78][12] = 1;dino_sprite[1][78][13] = 1;dino_sprite[1][78][14] = 1;dino_sprite[1][78][15] = 1;dino_sprite[1][78][16] = 1;dino_sprite[1][78][17] = 1;dino_sprite[1][78][18] = 1;dino_sprite[1][78][19] = 1;dino_sprite[1][78][20] = 1;dino_sprite[1][78][21] = 1;dino_sprite[1][78][22] = 1;dino_sprite[1][78][23] = 1;dino_sprite[1][78][24] = 1;dino_sprite[1][78][25] = 1;dino_sprite[1][78][29] = 1;dino_sprite[1][78][30] = 1;dino_sprite[1][78][31] = 1;dino_sprite[1][78][32] = 1;dino_sprite[1][78][33] = 1;dino_sprite[1][78][34] = 1;dino_sprite[1][78][35] = 1;dino_sprite[1][78][43] = 1;dino_sprite[1][78][44] = 1;dino_sprite[1][78][45] = 1;dino_sprite[1][78][46] = 1;dino_sprite[1][78][47] = 1;dino_sprite[1][78][48] = 1;dino_sprite[1][78][49] = 1;dino_sprite[1][78][50] = 1;dino_sprite[1][78][51] = 1;dino_sprite[1][78][52] = 1;dino_sprite[1][78][53] = 1;dino_sprite[1][78][54] = 1;dino_sprite[1][79][0] = 1;dino_sprite[1][79][1] = 1;dino_sprite[1][79][2] = 1;dino_sprite[1][79][3] = 1;dino_sprite[1][79][4] = 1;dino_sprite[1][79][5] = 1;dino_sprite[1][79][6] = 1;dino_sprite[1][79][7] = 1;dino_sprite[1][79][8] = 1;dino_sprite[1][79][9] = 1;dino_sprite[1][79][10] = 1;dino_sprite[1][79][11] = 1;dino_sprite[1][79][12] = 1;dino_sprite[1][79][13] = 1;dino_sprite[1][79][14] = 1;dino_sprite[1][79][15] = 1;dino_sprite[1][79][16] = 1;dino_sprite[1][79][17] = 1;dino_sprite[1][79][18] = 1;dino_sprite[1][79][19] = 1;dino_sprite[1][79][20] = 1;dino_sprite[1][79][21] = 1;dino_sprite[1][79][22] = 1;dino_sprite[1][79][23] = 1;dino_sprite[1][79][24] = 1;dino_sprite[1][79][25] = 1;dino_sprite[1][79][29] = 1;dino_sprite[1][79][30] = 1;dino_sprite[1][79][31] = 1;dino_sprite[1][79][32] = 1;dino_sprite[1][79][33] = 1;dino_sprite[1][79][34] = 1;dino_sprite[1][79][35] = 1;dino_sprite[1][79][43] = 1;dino_sprite[1][79][44] = 1;dino_sprite[1][79][45] = 1;dino_sprite[1][79][46] = 1;dino_sprite[1][79][47] = 1;dino_sprite[1][79][48] = 1;dino_sprite[1][79][49] = 1;dino_sprite[1][79][50] = 1;dino_sprite[1][79][51] = 1;dino_sprite[1][79][52] = 1;dino_sprite[1][79][53] = 1;dino_sprite[1][79][54] = 1;dino_sprite[1][80][0] = 1;dino_sprite[1][80][1] = 1;dino_sprite[1][80][2] = 1;dino_sprite[1][80][3] = 1;dino_sprite[1][80][4] = 1;dino_sprite[1][80][5] = 1;dino_sprite[1][80][6] = 1;dino_sprite[1][80][7] = 1;dino_sprite[1][80][8] = 1;dino_sprite[1][80][9] = 1;dino_sprite[1][80][10] = 1;dino_sprite[1][80][11] = 1;dino_sprite[1][80][12] = 1;dino_sprite[1][80][13] = 1;dino_sprite[1][80][14] = 1;dino_sprite[1][80][15] = 1;dino_sprite[1][80][16] = 1;dino_sprite[1][80][17] = 1;dino_sprite[1][80][18] = 1;dino_sprite[1][80][19] = 1;dino_sprite[1][80][20] = 1;dino_sprite[1][80][21] = 1;dino_sprite[1][80][22] = 1;dino_sprite[1][80][23] = 1;dino_sprite[1][80][24] = 1;dino_sprite[1][80][25] = 1;dino_sprite[1][80][29] = 1;dino_sprite[1][80][30] = 1;dino_sprite[1][80][31] = 1;dino_sprite[1][80][32] = 1;dino_sprite[1][80][33] = 1;dino_sprite[1][80][34] = 1;dino_sprite[1][80][35] = 1;dino_sprite[1][80][43] = 1;dino_sprite[1][80][44] = 1;dino_sprite[1][80][45] = 1;dino_sprite[1][80][46] = 1;dino_sprite[1][80][47] = 1;dino_sprite[1][80][48] = 1;dino_sprite[1][80][49] = 1;dino_sprite[1][80][50] = 1;dino_sprite[1][80][51] = 1;dino_sprite[1][80][52] = 1;dino_sprite[1][80][53] = 1;dino_sprite[1][80][54] = 1;dino_sprite[1][81][0] = 1;dino_sprite[1][81][1] = 1;dino_sprite[1][81][2] = 1;dino_sprite[1][81][3] = 1;dino_sprite[1][81][4] = 1;dino_sprite[1][81][5] = 1;dino_sprite[1][81][6] = 1;dino_sprite[1][81][7] = 1;dino_sprite[1][81][8] = 1;dino_sprite[1][81][9] = 1;dino_sprite[1][81][10] = 1;dino_sprite[1][81][11] = 1;dino_sprite[1][81][12] = 1;dino_sprite[1][81][13] = 1;dino_sprite[1][81][14] = 1;dino_sprite[1][81][15] = 1;dino_sprite[1][81][16] = 1;dino_sprite[1][81][17] = 1;dino_sprite[1][81][18] = 1;dino_sprite[1][81][19] = 1;dino_sprite[1][81][20] = 1;dino_sprite[1][81][21] = 1;dino_sprite[1][81][22] = 1;dino_sprite[1][81][23] = 1;dino_sprite[1][81][24] = 1;dino_sprite[1][81][25] = 1;dino_sprite[1][81][29] = 1;dino_sprite[1][81][30] = 1;dino_sprite[1][81][31] = 1;dino_sprite[1][81][32] = 1;dino_sprite[1][81][33] = 1;dino_sprite[1][81][34] = 1;dino_sprite[1][81][35] = 1;dino_sprite[1][81][43] = 1;dino_sprite[1][81][44] = 1;dino_sprite[1][81][45] = 1;dino_sprite[1][81][46] = 1;dino_sprite[1][81][47] = 1;dino_sprite[1][81][48] = 1;dino_sprite[1][81][49] = 1;dino_sprite[1][81][50] = 1;dino_sprite[1][81][51] = 1;dino_sprite[1][81][52] = 1;dino_sprite[1][81][53] = 1;dino_sprite[1][81][54] = 1;dino_sprite[1][82][0] = 1;dino_sprite[1][82][1] = 1;dino_sprite[1][82][2] = 1;dino_sprite[1][82][3] = 1;dino_sprite[1][82][4] = 1;dino_sprite[1][82][5] = 1;dino_sprite[1][82][6] = 1;dino_sprite[1][82][7] = 1;dino_sprite[1][82][8] = 1;dino_sprite[1][82][9] = 1;dino_sprite[1][82][10] = 1;dino_sprite[1][82][11] = 1;dino_sprite[1][82][12] = 1;dino_sprite[1][82][13] = 1;dino_sprite[1][82][14] = 1;dino_sprite[1][82][15] = 1;dino_sprite[1][82][16] = 1;dino_sprite[1][82][17] = 1;dino_sprite[1][82][18] = 1;dino_sprite[1][82][19] = 1;dino_sprite[1][82][20] = 1;dino_sprite[1][82][21] = 1;dino_sprite[1][82][22] = 1;dino_sprite[1][82][23] = 1;dino_sprite[1][82][24] = 1;dino_sprite[1][82][25] = 1;dino_sprite[1][82][29] = 1;dino_sprite[1][82][30] = 1;dino_sprite[1][82][31] = 1;dino_sprite[1][82][32] = 1;dino_sprite[1][82][33] = 1;dino_sprite[1][82][34] = 1;dino_sprite[1][82][35] = 1;dino_sprite[1][83][0] = 1;dino_sprite[1][83][1] = 1;dino_sprite[1][83][2] = 1;dino_sprite[1][83][3] = 1;dino_sprite[1][83][4] = 1;dino_sprite[1][83][5] = 1;dino_sprite[1][83][6] = 1;dino_sprite[1][83][7] = 1;dino_sprite[1][83][8] = 1;dino_sprite[1][83][9] = 1;dino_sprite[1][83][10] = 1;dino_sprite[1][83][11] = 1;dino_sprite[1][83][12] = 1;dino_sprite[1][83][13] = 1;dino_sprite[1][83][14] = 1;dino_sprite[1][83][15] = 1;dino_sprite[1][83][16] = 1;dino_sprite[1][83][17] = 1;dino_sprite[1][83][18] = 1;dino_sprite[1][83][19] = 1;dino_sprite[1][83][20] = 1;dino_sprite[1][83][21] = 1;dino_sprite[1][83][22] = 1;dino_sprite[1][83][23] = 1;dino_sprite[1][83][24] = 1;dino_sprite[1][83][25] = 1;dino_sprite[1][83][29] = 1;dino_sprite[1][83][30] = 1;dino_sprite[1][83][31] = 1;dino_sprite[1][83][32] = 1;dino_sprite[1][83][33] = 1;dino_sprite[1][83][34] = 1;dino_sprite[1][83][35] = 1;dino_sprite[1][84][0] = 1;dino_sprite[1][84][1] = 1;dino_sprite[1][84][2] = 1;dino_sprite[1][84][3] = 1;dino_sprite[1][84][4] = 1;dino_sprite[1][84][5] = 1;dino_sprite[1][84][6] = 1;dino_sprite[1][84][7] = 1;dino_sprite[1][84][8] = 1;dino_sprite[1][84][9] = 1;dino_sprite[1][84][10] = 1;dino_sprite[1][84][11] = 1;dino_sprite[1][84][12] = 1;dino_sprite[1][84][13] = 1;dino_sprite[1][84][14] = 1;dino_sprite[1][84][15] = 1;dino_sprite[1][84][16] = 1;dino_sprite[1][84][17] = 1;dino_sprite[1][84][18] = 1;dino_sprite[1][84][19] = 1;dino_sprite[1][84][20] = 1;dino_sprite[1][84][21] = 1;dino_sprite[1][84][22] = 1;dino_sprite[1][84][23] = 1;dino_sprite[1][84][24] = 1;dino_sprite[1][84][25] = 1;dino_sprite[1][84][29] = 1;dino_sprite[1][84][30] = 1;dino_sprite[1][84][31] = 1;dino_sprite[1][84][32] = 1;dino_sprite[1][84][33] = 1;dino_sprite[1][84][34] = 1;dino_sprite[1][84][35] = 1;dino_sprite[1][85][0] = 1;dino_sprite[1][85][1] = 1;dino_sprite[1][85][2] = 1;dino_sprite[1][85][3] = 1;dino_sprite[1][85][4] = 1;dino_sprite[1][85][5] = 1;dino_sprite[1][85][6] = 1;dino_sprite[1][85][7] = 1;dino_sprite[1][85][8] = 1;dino_sprite[1][85][9] = 1;dino_sprite[1][85][10] = 1;dino_sprite[1][85][11] = 1;dino_sprite[1][85][12] = 1;dino_sprite[1][85][13] = 1;dino_sprite[1][85][14] = 1;dino_sprite[1][85][15] = 1;dino_sprite[1][85][16] = 1;dino_sprite[1][85][17] = 1;dino_sprite[1][85][18] = 1;dino_sprite[1][85][19] = 1;dino_sprite[1][85][20] = 1;dino_sprite[1][85][21] = 1;dino_sprite[1][85][22] = 1;dino_sprite[1][85][23] = 1;dino_sprite[1][85][24] = 1;dino_sprite[1][85][25] = 1;dino_sprite[1][85][29] = 1;dino_sprite[1][85][30] = 1;dino_sprite[1][85][31] = 1;dino_sprite[1][85][32] = 1;dino_sprite[1][85][33] = 1;dino_sprite[1][85][34] = 1;dino_sprite[1][85][35] = 1;dino_sprite[1][86][0] = 1;dino_sprite[1][86][1] = 1;dino_sprite[1][86][2] = 1;dino_sprite[1][86][3] = 1;dino_sprite[1][86][4] = 1;dino_sprite[1][86][5] = 1;dino_sprite[1][86][6] = 1;dino_sprite[1][86][7] = 1;dino_sprite[1][86][8] = 1;dino_sprite[1][86][9] = 1;dino_sprite[1][86][10] = 1;dino_sprite[1][86][11] = 1;dino_sprite[1][86][12] = 1;dino_sprite[1][86][13] = 1;dino_sprite[1][86][14] = 1;dino_sprite[1][86][15] = 1;dino_sprite[1][86][16] = 1;dino_sprite[1][86][17] = 1;dino_sprite[1][86][18] = 1;dino_sprite[1][86][19] = 1;dino_sprite[1][86][20] = 1;dino_sprite[1][86][21] = 1;dino_sprite[1][86][22] = 1;dino_sprite[1][86][23] = 1;dino_sprite[1][86][24] = 1;dino_sprite[1][86][25] = 1;dino_sprite[1][86][29] = 1;dino_sprite[1][86][30] = 1;dino_sprite[1][86][31] = 1;dino_sprite[1][86][32] = 1;dino_sprite[1][86][33] = 1;dino_sprite[1][86][34] = 1;dino_sprite[1][86][35] = 1;dino_sprite[1][87][0] = 1;dino_sprite[1][87][1] = 1;dino_sprite[1][87][2] = 1;dino_sprite[1][87][3] = 1;dino_sprite[1][87][4] = 1;dino_sprite[1][87][5] = 1;dino_sprite[1][87][6] = 1;dino_sprite[1][87][7] = 1;dino_sprite[1][87][8] = 1;dino_sprite[1][87][9] = 1;dino_sprite[1][87][10] = 1;dino_sprite[1][87][11] = 1;dino_sprite[1][87][12] = 1;dino_sprite[1][87][13] = 1;dino_sprite[1][87][14] = 1;dino_sprite[1][87][15] = 1;dino_sprite[1][87][16] = 1;dino_sprite[1][87][17] = 1;dino_sprite[1][87][18] = 1;dino_sprite[1][87][19] = 1;dino_sprite[1][87][20] = 1;dino_sprite[1][87][21] = 1;dino_sprite[1][87][22] = 1;dino_sprite[1][87][23] = 1;dino_sprite[1][87][24] = 1;dino_sprite[1][87][25] = 1;dino_sprite[1][87][29] = 1;dino_sprite[1][87][30] = 1;dino_sprite[1][87][31] = 1;dino_sprite[1][87][32] = 1;dino_sprite[1][87][33] = 1;dino_sprite[1][87][34] = 1;dino_sprite[1][87][35] = 1;dino_sprite[1][88][0] = 1;dino_sprite[1][88][1] = 1;dino_sprite[1][88][2] = 1;dino_sprite[1][88][3] = 1;dino_sprite[1][88][4] = 1;dino_sprite[1][88][5] = 1;dino_sprite[1][88][6] = 1;dino_sprite[1][88][7] = 1;dino_sprite[1][88][8] = 1;dino_sprite[1][88][9] = 1;dino_sprite[1][88][10] = 1;dino_sprite[1][88][11] = 1;dino_sprite[1][88][12] = 1;dino_sprite[1][88][13] = 1;dino_sprite[1][88][14] = 1;dino_sprite[1][88][15] = 1;dino_sprite[1][88][16] = 1;dino_sprite[1][88][17] = 1;dino_sprite[1][88][18] = 1;dino_sprite[1][88][19] = 1;dino_sprite[1][88][20] = 1;dino_sprite[1][88][21] = 1;dino_sprite[1][88][22] = 1;dino_sprite[1][88][23] = 1;dino_sprite[1][88][24] = 1;dino_sprite[1][88][25] = 1;dino_sprite[1][88][29] = 1;dino_sprite[1][88][30] = 1;dino_sprite[1][88][31] = 1;dino_sprite[1][88][32] = 1;dino_sprite[1][88][33] = 1;dino_sprite[1][88][34] = 1;dino_sprite[1][88][35] = 1;dino_sprite[1][89][0] = 1;dino_sprite[1][89][1] = 1;dino_sprite[1][89][2] = 1;dino_sprite[1][89][3] = 1;dino_sprite[1][89][4] = 1;dino_sprite[1][89][5] = 1;dino_sprite[1][89][6] = 1;dino_sprite[1][89][7] = 1;dino_sprite[1][89][8] = 1;dino_sprite[1][89][9] = 1;dino_sprite[1][89][10] = 1;dino_sprite[1][89][11] = 1;dino_sprite[1][89][12] = 1;dino_sprite[1][89][13] = 1;dino_sprite[1][89][14] = 1;dino_sprite[1][89][15] = 1;dino_sprite[1][89][16] = 1;dino_sprite[1][89][17] = 1;dino_sprite[1][89][18] = 1;dino_sprite[1][89][19] = 1;dino_sprite[1][89][20] = 1;dino_sprite[1][89][21] = 1;dino_sprite[1][89][22] = 1;dino_sprite[1][89][23] = 1;dino_sprite[1][89][24] = 1;dino_sprite[1][89][25] = 1;dino_sprite[1][89][29] = 1;dino_sprite[1][89][30] = 1;dino_sprite[1][89][31] = 1;dino_sprite[1][89][32] = 1;dino_sprite[1][89][33] = 1;dino_sprite[1][89][34] = 1;dino_sprite[1][89][35] = 1;dino_sprite[1][90][0] = 1;dino_sprite[1][90][1] = 1;dino_sprite[1][90][2] = 1;dino_sprite[1][90][3] = 1;dino_sprite[1][90][4] = 1;dino_sprite[1][90][5] = 1;dino_sprite[1][90][6] = 1;dino_sprite[1][90][7] = 1;dino_sprite[1][90][8] = 1;dino_sprite[1][90][9] = 1;dino_sprite[1][90][10] = 1;dino_sprite[1][90][11] = 1;dino_sprite[1][90][12] = 1;dino_sprite[1][90][13] = 1;dino_sprite[1][90][14] = 1;dino_sprite[1][90][15] = 1;dino_sprite[1][90][16] = 1;dino_sprite[1][90][17] = 1;dino_sprite[1][90][18] = 1;dino_sprite[1][90][19] = 1;dino_sprite[1][90][20] = 1;dino_sprite[1][90][21] = 1;dino_sprite[1][90][22] = 1;dino_sprite[1][90][23] = 1;dino_sprite[1][90][24] = 1;dino_sprite[1][90][25] = 1;dino_sprite[1][90][29] = 1;dino_sprite[1][90][30] = 1;dino_sprite[1][90][31] = 1;dino_sprite[1][90][32] = 1;dino_sprite[1][90][33] = 1;dino_sprite[1][90][34] = 1;dino_sprite[1][90][35] = 1;dino_sprite[1][91][0] = 1;dino_sprite[1][91][1] = 1;dino_sprite[1][91][2] = 1;dino_sprite[1][91][3] = 1;dino_sprite[1][91][4] = 1;dino_sprite[1][91][5] = 1;dino_sprite[1][91][6] = 1;dino_sprite[1][91][7] = 1;dino_sprite[1][91][8] = 1;dino_sprite[1][91][9] = 1;dino_sprite[1][91][10] = 1;dino_sprite[1][91][11] = 1;dino_sprite[1][91][12] = 1;dino_sprite[1][91][13] = 1;dino_sprite[1][91][14] = 1;dino_sprite[1][91][15] = 1;dino_sprite[1][91][16] = 1;dino_sprite[1][91][17] = 1;dino_sprite[1][91][18] = 1;dino_sprite[1][91][19] = 1;dino_sprite[1][91][20] = 1;dino_sprite[1][91][21] = 1;dino_sprite[1][91][22] = 1;dino_sprite[1][91][23] = 1;dino_sprite[1][91][24] = 1;dino_sprite[1][91][25] = 1;dino_sprite[1][91][30] = 1;dino_sprite[1][91][31] = 1;dino_sprite[1][91][32] = 1;dino_sprite[1][91][33] = 1;dino_sprite[1][92][0] = 1;dino_sprite[1][92][1] = 1;dino_sprite[1][92][2] = 1;dino_sprite[1][92][3] = 1;dino_sprite[1][92][4] = 1;dino_sprite[1][92][5] = 1;dino_sprite[1][92][6] = 1;dino_sprite[1][92][7] = 1;dino_sprite[1][92][8] = 1;dino_sprite[1][92][9] = 1;dino_sprite[1][92][10] = 1;dino_sprite[1][92][11] = 1;dino_sprite[1][92][12] = 1;dino_sprite[1][92][13] = 1;dino_sprite[1][92][14] = 1;dino_sprite[1][92][15] = 1;dino_sprite[1][92][16] = 1;dino_sprite[1][92][17] = 1;dino_sprite[1][92][18] = 1;dino_sprite[1][92][19] = 1;dino_sprite[1][92][20] = 1;dino_sprite[1][92][21] = 1;dino_sprite[1][92][22] = 1;dino_sprite[1][92][23] = 1;dino_sprite[1][92][24] = 1;dino_sprite[1][92][25] = 1;dino_sprite[1][93][0] = 1;dino_sprite[1][93][1] = 1;dino_sprite[1][93][2] = 1;dino_sprite[1][93][3] = 1;dino_sprite[1][93][4] = 1;dino_sprite[1][93][5] = 1;dino_sprite[1][93][6] = 1;dino_sprite[1][93][7] = 1;dino_sprite[1][93][8] = 1;dino_sprite[1][93][9] = 1;dino_sprite[1][93][10] = 1;dino_sprite[1][93][11] = 1;dino_sprite[1][93][12] = 1;dino_sprite[1][93][13] = 1;dino_sprite[1][93][14] = 1;dino_sprite[1][93][15] = 1;dino_sprite[1][93][16] = 1;dino_sprite[1][93][17] = 1;dino_sprite[1][93][18] = 1;dino_sprite[1][93][19] = 1;dino_sprite[1][93][20] = 1;dino_sprite[1][93][21] = 1;dino_sprite[1][93][22] = 1;dino_sprite[1][93][23] = 1;dino_sprite[1][93][24] = 1;dino_sprite[1][93][25] = 1;dino_sprite[1][94][0] = 1;dino_sprite[1][94][1] = 1;dino_sprite[1][94][2] = 1;dino_sprite[1][94][3] = 1;dino_sprite[1][94][4] = 1;dino_sprite[1][94][5] = 1;dino_sprite[1][94][6] = 1;dino_sprite[1][94][7] = 1;dino_sprite[1][94][8] = 1;dino_sprite[1][94][9] = 1;dino_sprite[1][94][10] = 1;dino_sprite[1][94][11] = 1;dino_sprite[1][94][12] = 1;dino_sprite[1][94][13] = 1;dino_sprite[1][94][14] = 1;dino_sprite[1][94][15] = 1;dino_sprite[1][94][16] = 1;dino_sprite[1][94][17] = 1;dino_sprite[1][94][18] = 1;dino_sprite[1][94][19] = 1;dino_sprite[1][94][20] = 1;dino_sprite[1][94][21] = 1;dino_sprite[1][94][22] = 1;dino_sprite[1][94][23] = 1;dino_sprite[1][94][24] = 1;dino_sprite[1][94][25] = 1;dino_sprite[1][95][0] = 1;dino_sprite[1][95][1] = 1;dino_sprite[1][95][2] = 1;dino_sprite[1][95][3] = 1;dino_sprite[1][95][4] = 1;dino_sprite[1][95][5] = 1;dino_sprite[1][95][6] = 1;dino_sprite[1][95][7] = 1;dino_sprite[1][95][8] = 1;dino_sprite[1][95][9] = 1;dino_sprite[1][95][10] = 1;dino_sprite[1][95][11] = 1;dino_sprite[1][95][12] = 1;dino_sprite[1][95][13] = 1;dino_sprite[1][95][14] = 1;dino_sprite[1][95][15] = 1;dino_sprite[1][95][16] = 1;dino_sprite[1][95][17] = 1;dino_sprite[1][95][18] = 1;dino_sprite[1][95][19] = 1;dino_sprite[1][95][20] = 1;dino_sprite[1][95][21] = 1;dino_sprite[1][95][22] = 1;dino_sprite[1][95][23] = 1;dino_sprite[1][95][24] = 1;dino_sprite[1][95][25] = 1;dino_sprite[1][96][3] = 1;dino_sprite[1][96][4] = 1;dino_sprite[1][96][5] = 1;dino_sprite[1][96][6] = 1;dino_sprite[1][96][7] = 1;dino_sprite[1][96][8] = 1;dino_sprite[1][96][9] = 1;dino_sprite[1][96][10] = 1;dino_sprite[1][96][11] = 1;dino_sprite[1][96][12] = 1;dino_sprite[1][96][13] = 1;dino_sprite[1][96][14] = 1;dino_sprite[1][96][15] = 1;dino_sprite[1][96][16] = 1;dino_sprite[1][96][17] = 1;dino_sprite[1][96][18] = 1;dino_sprite[1][96][19] = 1;dino_sprite[1][96][20] = 1;dino_sprite[1][96][21] = 1;dino_sprite[1][96][22] = 1;dino_sprite[1][96][23] = 1;dino_sprite[1][96][24] = 1;dino_sprite[1][96][25] = 1;dino_sprite[1][97][3] = 1;dino_sprite[1][97][4] = 1;dino_sprite[1][97][5] = 1;dino_sprite[1][97][6] = 1;dino_sprite[1][97][7] = 1;dino_sprite[1][97][8] = 1;dino_sprite[1][97][9] = 1;dino_sprite[1][97][10] = 1;dino_sprite[1][97][11] = 1;dino_sprite[1][97][12] = 1;dino_sprite[1][97][13] = 1;dino_sprite[1][97][14] = 1;dino_sprite[1][97][15] = 1;dino_sprite[1][97][16] = 1;dino_sprite[1][97][17] = 1;dino_sprite[1][97][18] = 1;dino_sprite[1][97][19] = 1;dino_sprite[1][97][20] = 1;dino_sprite[1][97][21] = 1;dino_sprite[1][97][22] = 1;dino_sprite[1][97][23] = 1;dino_sprite[1][97][24] = 1;dino_sprite[1][97][25] = 1;dino_sprite[1][98][3] = 1;dino_sprite[1][98][4] = 1;dino_sprite[1][98][5] = 1;dino_sprite[1][98][6] = 1;dino_sprite[1][98][7] = 1;dino_sprite[1][98][8] = 1;dino_sprite[1][98][9] = 1;dino_sprite[1][98][10] = 1;dino_sprite[1][98][11] = 1;dino_sprite[1][98][12] = 1;dino_sprite[1][98][13] = 1;dino_sprite[1][98][14] = 1;dino_sprite[1][98][15] = 1;dino_sprite[1][98][16] = 1;dino_sprite[1][98][17] = 1;dino_sprite[1][98][18] = 1;dino_sprite[1][98][19] = 1;dino_sprite[1][98][20] = 1;dino_sprite[1][98][21] = 1;dino_sprite[1][98][22] = 1;dino_sprite[1][98][23] = 1;dino_sprite[1][98][24] = 1;dino_sprite[1][98][25] = 1;
	dino_sprite[2][2][35] = 1;dino_sprite[2][2][36] = 1;dino_sprite[2][2][37] = 1;dino_sprite[2][2][38] = 1;dino_sprite[2][2][39] = 1;dino_sprite[2][2][40] = 1;dino_sprite[2][2][41] = 1;dino_sprite[2][2][42] = 1;dino_sprite[2][2][43] = 1;dino_sprite[2][2][44] = 1;dino_sprite[2][2][45] = 1;dino_sprite[2][2][46] = 1;dino_sprite[2][2][47] = 1;dino_sprite[2][2][48] = 1;dino_sprite[2][2][49] = 1;dino_sprite[2][2][50] = 1;dino_sprite[2][2][51] = 1;dino_sprite[2][2][52] = 1;dino_sprite[2][2][53] = 1;dino_sprite[2][2][54] = 1;dino_sprite[2][2][55] = 1;dino_sprite[2][2][56] = 1;dino_sprite[2][2][57] = 1;dino_sprite[2][2][58] = 1;dino_sprite[2][2][59] = 1;dino_sprite[2][2][60] = 1;dino_sprite[2][2][61] = 1;dino_sprite[2][2][62] = 1;dino_sprite[2][3][35] = 1;dino_sprite[2][3][36] = 1;dino_sprite[2][3][37] = 1;dino_sprite[2][3][38] = 1;dino_sprite[2][3][39] = 1;dino_sprite[2][3][40] = 1;dino_sprite[2][3][41] = 1;dino_sprite[2][3][42] = 1;dino_sprite[2][3][43] = 1;dino_sprite[2][3][44] = 1;dino_sprite[2][3][45] = 1;dino_sprite[2][3][46] = 1;dino_sprite[2][3][47] = 1;dino_sprite[2][3][48] = 1;dino_sprite[2][3][49] = 1;dino_sprite[2][3][50] = 1;dino_sprite[2][3][51] = 1;dino_sprite[2][3][52] = 1;dino_sprite[2][3][53] = 1;dino_sprite[2][3][54] = 1;dino_sprite[2][3][55] = 1;dino_sprite[2][3][56] = 1;dino_sprite[2][3][57] = 1;dino_sprite[2][3][58] = 1;dino_sprite[2][3][59] = 1;dino_sprite[2][3][60] = 1;dino_sprite[2][3][61] = 1;dino_sprite[2][3][62] = 1;dino_sprite[2][4][35] = 1;dino_sprite[2][4][36] = 1;dino_sprite[2][4][37] = 1;dino_sprite[2][4][38] = 1;dino_sprite[2][4][39] = 1;dino_sprite[2][4][40] = 1;dino_sprite[2][4][41] = 1;dino_sprite[2][4][42] = 1;dino_sprite[2][4][43] = 1;dino_sprite[2][4][44] = 1;dino_sprite[2][4][45] = 1;dino_sprite[2][4][46] = 1;dino_sprite[2][4][47] = 1;dino_sprite[2][4][48] = 1;dino_sprite[2][4][49] = 1;dino_sprite[2][4][50] = 1;dino_sprite[2][4][51] = 1;dino_sprite[2][4][52] = 1;dino_sprite[2][4][53] = 1;dino_sprite[2][4][54] = 1;dino_sprite[2][4][55] = 1;dino_sprite[2][4][56] = 1;dino_sprite[2][4][57] = 1;dino_sprite[2][4][58] = 1;dino_sprite[2][4][59] = 1;dino_sprite[2][4][60] = 1;dino_sprite[2][4][61] = 1;dino_sprite[2][4][62] = 1;dino_sprite[2][5][35] = 1;dino_sprite[2][5][36] = 1;dino_sprite[2][5][37] = 1;dino_sprite[2][5][38] = 1;dino_sprite[2][5][39] = 1;dino_sprite[2][5][40] = 1;dino_sprite[2][5][41] = 1;dino_sprite[2][5][42] = 1;dino_sprite[2][5][43] = 1;dino_sprite[2][5][44] = 1;dino_sprite[2][5][45] = 1;dino_sprite[2][5][46] = 1;dino_sprite[2][5][47] = 1;dino_sprite[2][5][48] = 1;dino_sprite[2][5][49] = 1;dino_sprite[2][5][50] = 1;dino_sprite[2][5][51] = 1;dino_sprite[2][5][52] = 1;dino_sprite[2][5][53] = 1;dino_sprite[2][5][54] = 1;dino_sprite[2][5][55] = 1;dino_sprite[2][5][56] = 1;dino_sprite[2][5][57] = 1;dino_sprite[2][5][58] = 1;dino_sprite[2][5][59] = 1;dino_sprite[2][5][60] = 1;dino_sprite[2][5][61] = 1;dino_sprite[2][5][62] = 1;dino_sprite[2][6][35] = 1;dino_sprite[2][6][36] = 1;dino_sprite[2][6][37] = 1;dino_sprite[2][6][38] = 1;dino_sprite[2][6][39] = 1;dino_sprite[2][6][40] = 1;dino_sprite[2][6][41] = 1;dino_sprite[2][6][42] = 1;dino_sprite[2][6][43] = 1;dino_sprite[2][6][44] = 1;dino_sprite[2][6][45] = 1;dino_sprite[2][6][46] = 1;dino_sprite[2][6][47] = 1;dino_sprite[2][6][48] = 1;dino_sprite[2][6][49] = 1;dino_sprite[2][6][50] = 1;dino_sprite[2][6][51] = 1;dino_sprite[2][6][52] = 1;dino_sprite[2][6][53] = 1;dino_sprite[2][6][54] = 1;dino_sprite[2][6][55] = 1;dino_sprite[2][6][56] = 1;dino_sprite[2][6][57] = 1;dino_sprite[2][6][58] = 1;dino_sprite[2][6][59] = 1;dino_sprite[2][6][60] = 1;dino_sprite[2][6][61] = 1;dino_sprite[2][6][62] = 1;dino_sprite[2][7][35] = 1;dino_sprite[2][7][36] = 1;dino_sprite[2][7][37] = 1;dino_sprite[2][7][38] = 1;dino_sprite[2][7][39] = 1;dino_sprite[2][7][40] = 1;dino_sprite[2][7][41] = 1;dino_sprite[2][7][42] = 1;dino_sprite[2][7][43] = 1;dino_sprite[2][7][44] = 1;dino_sprite[2][7][45] = 1;dino_sprite[2][7][46] = 1;dino_sprite[2][7][47] = 1;dino_sprite[2][7][48] = 1;dino_sprite[2][7][49] = 1;dino_sprite[2][7][50] = 1;dino_sprite[2][7][51] = 1;dino_sprite[2][7][52] = 1;dino_sprite[2][7][53] = 1;dino_sprite[2][7][54] = 1;dino_sprite[2][7][55] = 1;dino_sprite[2][7][56] = 1;dino_sprite[2][7][57] = 1;dino_sprite[2][7][58] = 1;dino_sprite[2][7][59] = 1;dino_sprite[2][7][60] = 1;dino_sprite[2][7][61] = 1;dino_sprite[2][7][62] = 1;dino_sprite[2][7][63] = 1;dino_sprite[2][7][64] = 1;dino_sprite[2][7][65] = 1;dino_sprite[2][7][66] = 1;dino_sprite[2][7][67] = 1;dino_sprite[2][8][44] = 1;dino_sprite[2][8][45] = 1;dino_sprite[2][8][46] = 1;dino_sprite[2][8][47] = 1;dino_sprite[2][8][48] = 1;dino_sprite[2][8][49] = 1;dino_sprite[2][8][50] = 1;dino_sprite[2][8][51] = 1;dino_sprite[2][8][52] = 1;dino_sprite[2][8][53] = 1;dino_sprite[2][8][54] = 1;dino_sprite[2][8][55] = 1;dino_sprite[2][8][56] = 1;dino_sprite[2][8][57] = 1;dino_sprite[2][8][58] = 1;dino_sprite[2][8][59] = 1;dino_sprite[2][8][60] = 1;dino_sprite[2][8][61] = 1;dino_sprite[2][8][62] = 1;dino_sprite[2][8][63] = 1;dino_sprite[2][8][64] = 1;dino_sprite[2][8][65] = 1;dino_sprite[2][8][66] = 1;dino_sprite[2][8][67] = 1;dino_sprite[2][9][44] = 1;dino_sprite[2][9][45] = 1;dino_sprite[2][9][46] = 1;dino_sprite[2][9][47] = 1;dino_sprite[2][9][48] = 1;dino_sprite[2][9][49] = 1;dino_sprite[2][9][50] = 1;dino_sprite[2][9][51] = 1;dino_sprite[2][9][52] = 1;dino_sprite[2][9][53] = 1;dino_sprite[2][9][54] = 1;dino_sprite[2][9][55] = 1;dino_sprite[2][9][56] = 1;dino_sprite[2][9][57] = 1;dino_sprite[2][9][58] = 1;dino_sprite[2][9][59] = 1;dino_sprite[2][9][60] = 1;dino_sprite[2][9][61] = 1;dino_sprite[2][9][62] = 1;dino_sprite[2][9][63] = 1;dino_sprite[2][9][64] = 1;dino_sprite[2][9][65] = 1;dino_sprite[2][9][66] = 1;dino_sprite[2][9][67] = 1;dino_sprite[2][10][44] = 1;dino_sprite[2][10][45] = 1;dino_sprite[2][10][46] = 1;dino_sprite[2][10][47] = 1;dino_sprite[2][10][48] = 1;dino_sprite[2][10][49] = 1;dino_sprite[2][10][50] = 1;dino_sprite[2][10][51] = 1;dino_sprite[2][10][52] = 1;dino_sprite[2][10][53] = 1;dino_sprite[2][10][54] = 1;dino_sprite[2][10][55] = 1;dino_sprite[2][10][56] = 1;dino_sprite[2][10][57] = 1;dino_sprite[2][10][58] = 1;dino_sprite[2][10][59] = 1;dino_sprite[2][10][60] = 1;dino_sprite[2][10][61] = 1;dino_sprite[2][10][62] = 1;dino_sprite[2][10][63] = 1;dino_sprite[2][10][64] = 1;dino_sprite[2][10][65] = 1;dino_sprite[2][10][66] = 1;dino_sprite[2][10][67] = 1;dino_sprite[2][11][44] = 1;dino_sprite[2][11][45] = 1;dino_sprite[2][11][46] = 1;dino_sprite[2][11][47] = 1;dino_sprite[2][11][48] = 1;dino_sprite[2][11][49] = 1;dino_sprite[2][11][50] = 1;dino_sprite[2][11][51] = 1;dino_sprite[2][11][52] = 1;dino_sprite[2][11][53] = 1;dino_sprite[2][11][54] = 1;dino_sprite[2][11][55] = 1;dino_sprite[2][11][56] = 1;dino_sprite[2][11][57] = 1;dino_sprite[2][11][58] = 1;dino_sprite[2][11][59] = 1;dino_sprite[2][11][60] = 1;dino_sprite[2][11][61] = 1;dino_sprite[2][11][62] = 1;dino_sprite[2][11][63] = 1;dino_sprite[2][11][64] = 1;dino_sprite[2][11][65] = 1;dino_sprite[2][11][66] = 1;dino_sprite[2][11][67] = 1;dino_sprite[2][12][49] = 1;dino_sprite[2][12][50] = 1;dino_sprite[2][12][51] = 1;dino_sprite[2][12][52] = 1;dino_sprite[2][12][53] = 1;dino_sprite[2][12][54] = 1;dino_sprite[2][12][55] = 1;dino_sprite[2][12][56] = 1;dino_sprite[2][12][57] = 1;dino_sprite[2][12][58] = 1;dino_sprite[2][12][59] = 1;dino_sprite[2][12][60] = 1;dino_sprite[2][12][61] = 1;dino_sprite[2][12][62] = 1;dino_sprite[2][12][63] = 1;dino_sprite[2][12][64] = 1;dino_sprite[2][12][65] = 1;dino_sprite[2][12][66] = 1;dino_sprite[2][12][67] = 1;dino_sprite[2][12][68] = 1;dino_sprite[2][12][69] = 1;dino_sprite[2][12][70] = 1;dino_sprite[2][12][71] = 1;dino_sprite[2][12][72] = 1;dino_sprite[2][13][49] = 1;dino_sprite[2][13][50] = 1;dino_sprite[2][13][51] = 1;dino_sprite[2][13][52] = 1;dino_sprite[2][13][53] = 1;dino_sprite[2][13][54] = 1;dino_sprite[2][13][55] = 1;dino_sprite[2][13][56] = 1;dino_sprite[2][13][57] = 1;dino_sprite[2][13][58] = 1;dino_sprite[2][13][59] = 1;dino_sprite[2][13][60] = 1;dino_sprite[2][13][61] = 1;dino_sprite[2][13][62] = 1;dino_sprite[2][13][63] = 1;dino_sprite[2][13][64] = 1;dino_sprite[2][13][65] = 1;dino_sprite[2][13][66] = 1;dino_sprite[2][13][67] = 1;dino_sprite[2][13][68] = 1;dino_sprite[2][13][69] = 1;dino_sprite[2][13][70] = 1;dino_sprite[2][13][71] = 1;dino_sprite[2][13][72] = 1;dino_sprite[2][14][49] = 1;dino_sprite[2][14][50] = 1;dino_sprite[2][14][51] = 1;dino_sprite[2][14][52] = 1;dino_sprite[2][14][53] = 1;dino_sprite[2][14][54] = 1;dino_sprite[2][14][55] = 1;dino_sprite[2][14][56] = 1;dino_sprite[2][14][57] = 1;dino_sprite[2][14][58] = 1;dino_sprite[2][14][59] = 1;dino_sprite[2][14][60] = 1;dino_sprite[2][14][61] = 1;dino_sprite[2][14][62] = 1;dino_sprite[2][14][63] = 1;dino_sprite[2][14][64] = 1;dino_sprite[2][14][65] = 1;dino_sprite[2][14][66] = 1;dino_sprite[2][14][67] = 1;dino_sprite[2][14][68] = 1;dino_sprite[2][14][69] = 1;dino_sprite[2][14][70] = 1;dino_sprite[2][14][71] = 1;dino_sprite[2][14][72] = 1;dino_sprite[2][15][49] = 1;dino_sprite[2][15][50] = 1;dino_sprite[2][15][51] = 1;dino_sprite[2][15][52] = 1;dino_sprite[2][15][53] = 1;dino_sprite[2][15][54] = 1;dino_sprite[2][15][55] = 1;dino_sprite[2][15][56] = 1;dino_sprite[2][15][57] = 1;dino_sprite[2][15][58] = 1;dino_sprite[2][15][59] = 1;dino_sprite[2][15][60] = 1;dino_sprite[2][15][61] = 1;dino_sprite[2][15][62] = 1;dino_sprite[2][15][63] = 1;dino_sprite[2][15][64] = 1;dino_sprite[2][15][65] = 1;dino_sprite[2][15][66] = 1;dino_sprite[2][15][67] = 1;dino_sprite[2][15][68] = 1;dino_sprite[2][15][69] = 1;dino_sprite[2][15][70] = 1;dino_sprite[2][15][71] = 1;dino_sprite[2][15][72] = 1;dino_sprite[2][16][49] = 1;dino_sprite[2][16][50] = 1;dino_sprite[2][16][51] = 1;dino_sprite[2][16][52] = 1;dino_sprite[2][16][53] = 1;dino_sprite[2][16][54] = 1;dino_sprite[2][16][55] = 1;dino_sprite[2][16][56] = 1;dino_sprite[2][16][57] = 1;dino_sprite[2][16][58] = 1;dino_sprite[2][16][59] = 1;dino_sprite[2][16][60] = 1;dino_sprite[2][16][61] = 1;dino_sprite[2][16][62] = 1;dino_sprite[2][16][63] = 1;dino_sprite[2][16][64] = 1;dino_sprite[2][16][65] = 1;dino_sprite[2][16][66] = 1;dino_sprite[2][16][67] = 1;dino_sprite[2][16][68] = 1;dino_sprite[2][16][69] = 1;dino_sprite[2][16][70] = 1;dino_sprite[2][16][71] = 1;dino_sprite[2][16][72] = 1;dino_sprite[2][17][54] = 1;dino_sprite[2][17][55] = 1;dino_sprite[2][17][56] = 1;dino_sprite[2][17][57] = 1;dino_sprite[2][17][58] = 1;dino_sprite[2][17][59] = 1;dino_sprite[2][17][60] = 1;dino_sprite[2][17][61] = 1;dino_sprite[2][17][62] = 1;dino_sprite[2][17][63] = 1;dino_sprite[2][17][64] = 1;dino_sprite[2][17][65] = 1;dino_sprite[2][17][66] = 1;dino_sprite[2][17][67] = 1;dino_sprite[2][17][68] = 1;dino_sprite[2][17][69] = 1;dino_sprite[2][17][70] = 1;dino_sprite[2][17][71] = 1;dino_sprite[2][17][72] = 1;dino_sprite[2][17][73] = 1;dino_sprite[2][17][74] = 1;dino_sprite[2][17][75] = 1;dino_sprite[2][17][76] = 1;dino_sprite[2][17][77] = 1;dino_sprite[2][18][54] = 1;dino_sprite[2][18][55] = 1;dino_sprite[2][18][56] = 1;dino_sprite[2][18][57] = 1;dino_sprite[2][18][58] = 1;dino_sprite[2][18][59] = 1;dino_sprite[2][18][60] = 1;dino_sprite[2][18][61] = 1;dino_sprite[2][18][62] = 1;dino_sprite[2][18][63] = 1;dino_sprite[2][18][64] = 1;dino_sprite[2][18][65] = 1;dino_sprite[2][18][66] = 1;dino_sprite[2][18][67] = 1;dino_sprite[2][18][68] = 1;dino_sprite[2][18][69] = 1;dino_sprite[2][18][70] = 1;dino_sprite[2][18][71] = 1;dino_sprite[2][18][72] = 1;dino_sprite[2][18][73] = 1;dino_sprite[2][18][74] = 1;dino_sprite[2][18][75] = 1;dino_sprite[2][18][76] = 1;dino_sprite[2][18][77] = 1;dino_sprite[2][19][54] = 1;dino_sprite[2][19][55] = 1;dino_sprite[2][19][56] = 1;dino_sprite[2][19][57] = 1;dino_sprite[2][19][58] = 1;dino_sprite[2][19][59] = 1;dino_sprite[2][19][60] = 1;dino_sprite[2][19][61] = 1;dino_sprite[2][19][62] = 1;dino_sprite[2][19][63] = 1;dino_sprite[2][19][64] = 1;dino_sprite[2][19][65] = 1;dino_sprite[2][19][66] = 1;dino_sprite[2][19][67] = 1;dino_sprite[2][19][68] = 1;dino_sprite[2][19][69] = 1;dino_sprite[2][19][70] = 1;dino_sprite[2][19][71] = 1;dino_sprite[2][19][72] = 1;dino_sprite[2][19][73] = 1;dino_sprite[2][19][74] = 1;dino_sprite[2][19][75] = 1;dino_sprite[2][19][76] = 1;dino_sprite[2][19][77] = 1;dino_sprite[2][20][54] = 1;dino_sprite[2][20][55] = 1;dino_sprite[2][20][56] = 1;dino_sprite[2][20][57] = 1;dino_sprite[2][20][58] = 1;dino_sprite[2][20][59] = 1;dino_sprite[2][20][60] = 1;dino_sprite[2][20][61] = 1;dino_sprite[2][20][62] = 1;dino_sprite[2][20][63] = 1;dino_sprite[2][20][64] = 1;dino_sprite[2][20][65] = 1;dino_sprite[2][20][66] = 1;dino_sprite[2][20][67] = 1;dino_sprite[2][20][68] = 1;dino_sprite[2][20][69] = 1;dino_sprite[2][20][70] = 1;dino_sprite[2][20][71] = 1;dino_sprite[2][20][72] = 1;dino_sprite[2][20][73] = 1;dino_sprite[2][20][74] = 1;dino_sprite[2][20][75] = 1;dino_sprite[2][20][76] = 1;dino_sprite[2][20][77] = 1;dino_sprite[2][21][54] = 1;dino_sprite[2][21][55] = 1;dino_sprite[2][21][56] = 1;dino_sprite[2][21][57] = 1;dino_sprite[2][21][58] = 1;dino_sprite[2][21][59] = 1;dino_sprite[2][21][60] = 1;dino_sprite[2][21][61] = 1;dino_sprite[2][21][62] = 1;dino_sprite[2][21][63] = 1;dino_sprite[2][21][64] = 1;dino_sprite[2][21][65] = 1;dino_sprite[2][21][66] = 1;dino_sprite[2][21][67] = 1;dino_sprite[2][21][68] = 1;dino_sprite[2][21][69] = 1;dino_sprite[2][21][70] = 1;dino_sprite[2][21][71] = 1;dino_sprite[2][21][72] = 1;dino_sprite[2][21][73] = 1;dino_sprite[2][21][74] = 1;dino_sprite[2][21][75] = 1;dino_sprite[2][21][76] = 1;dino_sprite[2][21][77] = 1;dino_sprite[2][22][54] = 1;dino_sprite[2][22][55] = 1;dino_sprite[2][22][56] = 1;dino_sprite[2][22][57] = 1;dino_sprite[2][22][58] = 1;dino_sprite[2][22][59] = 1;dino_sprite[2][22][60] = 1;dino_sprite[2][22][61] = 1;dino_sprite[2][22][62] = 1;dino_sprite[2][22][63] = 1;dino_sprite[2][22][64] = 1;dino_sprite[2][22][65] = 1;dino_sprite[2][22][66] = 1;dino_sprite[2][22][67] = 1;dino_sprite[2][22][68] = 1;dino_sprite[2][22][69] = 1;dino_sprite[2][22][70] = 1;dino_sprite[2][22][71] = 1;dino_sprite[2][22][72] = 1;dino_sprite[2][22][73] = 1;dino_sprite[2][22][74] = 1;dino_sprite[2][22][75] = 1;dino_sprite[2][22][76] = 1;dino_sprite[2][22][77] = 1;dino_sprite[2][22][78] = 1;dino_sprite[2][22][79] = 1;dino_sprite[2][22][80] = 1;dino_sprite[2][22][81] = 1;dino_sprite[2][23][54] = 1;dino_sprite[2][23][55] = 1;dino_sprite[2][23][56] = 1;dino_sprite[2][23][57] = 1;dino_sprite[2][23][58] = 1;dino_sprite[2][23][59] = 1;dino_sprite[2][23][60] = 1;dino_sprite[2][23][61] = 1;dino_sprite[2][23][62] = 1;dino_sprite[2][23][63] = 1;dino_sprite[2][23][64] = 1;dino_sprite[2][23][65] = 1;dino_sprite[2][23][66] = 1;dino_sprite[2][23][67] = 1;dino_sprite[2][23][68] = 1;dino_sprite[2][23][69] = 1;dino_sprite[2][23][70] = 1;dino_sprite[2][23][71] = 1;dino_sprite[2][23][72] = 1;dino_sprite[2][23][73] = 1;dino_sprite[2][23][74] = 1;dino_sprite[2][23][75] = 1;dino_sprite[2][23][76] = 1;dino_sprite[2][23][77] = 1;dino_sprite[2][23][78] = 1;dino_sprite[2][23][79] = 1;dino_sprite[2][23][80] = 1;dino_sprite[2][23][81] = 1;dino_sprite[2][24][54] = 1;dino_sprite[2][24][55] = 1;dino_sprite[2][24][56] = 1;dino_sprite[2][24][57] = 1;dino_sprite[2][24][58] = 1;dino_sprite[2][24][59] = 1;dino_sprite[2][24][60] = 1;dino_sprite[2][24][61] = 1;dino_sprite[2][24][62] = 1;dino_sprite[2][24][63] = 1;dino_sprite[2][24][64] = 1;dino_sprite[2][24][65] = 1;dino_sprite[2][24][66] = 1;dino_sprite[2][24][67] = 1;dino_sprite[2][24][68] = 1;dino_sprite[2][24][69] = 1;dino_sprite[2][24][70] = 1;dino_sprite[2][24][71] = 1;dino_sprite[2][24][72] = 1;dino_sprite[2][24][73] = 1;dino_sprite[2][24][74] = 1;dino_sprite[2][24][75] = 1;dino_sprite[2][24][76] = 1;dino_sprite[2][24][77] = 1;dino_sprite[2][24][78] = 1;dino_sprite[2][24][79] = 1;dino_sprite[2][24][80] = 1;dino_sprite[2][24][81] = 1;dino_sprite[2][25][54] = 1;dino_sprite[2][25][55] = 1;dino_sprite[2][25][56] = 1;dino_sprite[2][25][57] = 1;dino_sprite[2][25][58] = 1;dino_sprite[2][25][59] = 1;dino_sprite[2][25][60] = 1;dino_sprite[2][25][61] = 1;dino_sprite[2][25][62] = 1;dino_sprite[2][25][63] = 1;dino_sprite[2][25][64] = 1;dino_sprite[2][25][65] = 1;dino_sprite[2][25][66] = 1;dino_sprite[2][25][67] = 1;dino_sprite[2][25][68] = 1;dino_sprite[2][25][69] = 1;dino_sprite[2][25][70] = 1;dino_sprite[2][25][71] = 1;dino_sprite[2][25][72] = 1;dino_sprite[2][25][73] = 1;dino_sprite[2][25][74] = 1;dino_sprite[2][25][75] = 1;dino_sprite[2][25][76] = 1;dino_sprite[2][25][77] = 1;dino_sprite[2][25][78] = 1;dino_sprite[2][25][79] = 1;dino_sprite[2][25][80] = 1;dino_sprite[2][25][81] = 1;dino_sprite[2][26][49] = 1;dino_sprite[2][26][50] = 1;dino_sprite[2][26][51] = 1;dino_sprite[2][26][52] = 1;dino_sprite[2][26][53] = 1;dino_sprite[2][26][54] = 1;dino_sprite[2][26][55] = 1;dino_sprite[2][26][56] = 1;dino_sprite[2][26][57] = 1;dino_sprite[2][26][58] = 1;dino_sprite[2][26][59] = 1;dino_sprite[2][26][60] = 1;dino_sprite[2][26][61] = 1;dino_sprite[2][26][62] = 1;dino_sprite[2][26][63] = 1;dino_sprite[2][26][64] = 1;dino_sprite[2][26][65] = 1;dino_sprite[2][26][66] = 1;dino_sprite[2][26][67] = 1;dino_sprite[2][26][68] = 1;dino_sprite[2][26][69] = 1;dino_sprite[2][26][70] = 1;dino_sprite[2][26][71] = 1;dino_sprite[2][26][72] = 1;dino_sprite[2][26][73] = 1;dino_sprite[2][26][74] = 1;dino_sprite[2][26][75] = 1;dino_sprite[2][26][76] = 1;dino_sprite[2][26][77] = 1;dino_sprite[2][26][78] = 1;dino_sprite[2][26][79] = 1;dino_sprite[2][26][80] = 1;dino_sprite[2][26][81] = 1;dino_sprite[2][26][82] = 1;dino_sprite[2][26][83] = 1;dino_sprite[2][26][84] = 1;dino_sprite[2][26][85] = 1;dino_sprite[2][26][86] = 1;dino_sprite[2][26][87] = 1;dino_sprite[2][26][88] = 1;dino_sprite[2][26][89] = 1;dino_sprite[2][26][90] = 1;dino_sprite[2][26][91] = 1;dino_sprite[2][26][92] = 1;dino_sprite[2][26][93] = 1;dino_sprite[2][26][94] = 1;dino_sprite[2][26][95] = 1;dino_sprite[2][26][96] = 1;dino_sprite[2][26][97] = 1;dino_sprite[2][26][98] = 1;dino_sprite[2][26][99] = 1;dino_sprite[2][27][49] = 1;dino_sprite[2][27][50] = 1;dino_sprite[2][27][51] = 1;dino_sprite[2][27][52] = 1;dino_sprite[2][27][53] = 1;dino_sprite[2][27][54] = 1;dino_sprite[2][27][55] = 1;dino_sprite[2][27][56] = 1;dino_sprite[2][27][57] = 1;dino_sprite[2][27][58] = 1;dino_sprite[2][27][59] = 1;dino_sprite[2][27][60] = 1;dino_sprite[2][27][61] = 1;dino_sprite[2][27][62] = 1;dino_sprite[2][27][63] = 1;dino_sprite[2][27][64] = 1;dino_sprite[2][27][65] = 1;dino_sprite[2][27][66] = 1;dino_sprite[2][27][67] = 1;dino_sprite[2][27][68] = 1;dino_sprite[2][27][69] = 1;dino_sprite[2][27][70] = 1;dino_sprite[2][27][71] = 1;dino_sprite[2][27][72] = 1;dino_sprite[2][27][73] = 1;dino_sprite[2][27][74] = 1;dino_sprite[2][27][75] = 1;dino_sprite[2][27][76] = 1;dino_sprite[2][27][77] = 1;dino_sprite[2][27][78] = 1;dino_sprite[2][27][79] = 1;dino_sprite[2][27][80] = 1;dino_sprite[2][27][81] = 1;dino_sprite[2][27][82] = 1;dino_sprite[2][27][83] = 1;dino_sprite[2][27][84] = 1;dino_sprite[2][27][85] = 1;dino_sprite[2][27][86] = 1;dino_sprite[2][27][87] = 1;dino_sprite[2][27][88] = 1;dino_sprite[2][27][89] = 1;dino_sprite[2][27][90] = 1;dino_sprite[2][27][91] = 1;dino_sprite[2][27][92] = 1;dino_sprite[2][27][93] = 1;dino_sprite[2][27][94] = 1;dino_sprite[2][27][95] = 1;dino_sprite[2][27][96] = 1;dino_sprite[2][27][97] = 1;dino_sprite[2][27][98] = 1;dino_sprite[2][27][99] = 1;dino_sprite[2][28][49] = 1;dino_sprite[2][28][50] = 1;dino_sprite[2][28][51] = 1;dino_sprite[2][28][52] = 1;dino_sprite[2][28][53] = 1;dino_sprite[2][28][54] = 1;dino_sprite[2][28][55] = 1;dino_sprite[2][28][56] = 1;dino_sprite[2][28][57] = 1;dino_sprite[2][28][58] = 1;dino_sprite[2][28][59] = 1;dino_sprite[2][28][60] = 1;dino_sprite[2][28][61] = 1;dino_sprite[2][28][62] = 1;dino_sprite[2][28][63] = 1;dino_sprite[2][28][64] = 1;dino_sprite[2][28][65] = 1;dino_sprite[2][28][66] = 1;dino_sprite[2][28][67] = 1;dino_sprite[2][28][68] = 1;dino_sprite[2][28][69] = 1;dino_sprite[2][28][70] = 1;dino_sprite[2][28][71] = 1;dino_sprite[2][28][72] = 1;dino_sprite[2][28][73] = 1;dino_sprite[2][28][74] = 1;dino_sprite[2][28][75] = 1;dino_sprite[2][28][76] = 1;dino_sprite[2][28][77] = 1;dino_sprite[2][28][78] = 1;dino_sprite[2][28][79] = 1;dino_sprite[2][28][80] = 1;dino_sprite[2][28][81] = 1;dino_sprite[2][28][82] = 1;dino_sprite[2][28][83] = 1;dino_sprite[2][28][84] = 1;dino_sprite[2][28][85] = 1;dino_sprite[2][28][86] = 1;dino_sprite[2][28][87] = 1;dino_sprite[2][28][88] = 1;dino_sprite[2][28][89] = 1;dino_sprite[2][28][90] = 1;dino_sprite[2][28][91] = 1;dino_sprite[2][28][92] = 1;dino_sprite[2][28][93] = 1;dino_sprite[2][28][94] = 1;dino_sprite[2][28][95] = 1;dino_sprite[2][28][96] = 1;dino_sprite[2][28][97] = 1;dino_sprite[2][28][98] = 1;dino_sprite[2][28][99] = 1;dino_sprite[2][29][49] = 1;dino_sprite[2][29][50] = 1;dino_sprite[2][29][51] = 1;dino_sprite[2][29][52] = 1;dino_sprite[2][29][53] = 1;dino_sprite[2][29][54] = 1;dino_sprite[2][29][55] = 1;dino_sprite[2][29][56] = 1;dino_sprite[2][29][57] = 1;dino_sprite[2][29][58] = 1;dino_sprite[2][29][59] = 1;dino_sprite[2][29][60] = 1;dino_sprite[2][29][61] = 1;dino_sprite[2][29][62] = 1;dino_sprite[2][29][63] = 1;dino_sprite[2][29][64] = 1;dino_sprite[2][29][65] = 1;dino_sprite[2][29][66] = 1;dino_sprite[2][29][67] = 1;dino_sprite[2][29][68] = 1;dino_sprite[2][29][69] = 1;dino_sprite[2][29][70] = 1;dino_sprite[2][29][71] = 1;dino_sprite[2][29][72] = 1;dino_sprite[2][29][73] = 1;dino_sprite[2][29][74] = 1;dino_sprite[2][29][75] = 1;dino_sprite[2][29][76] = 1;dino_sprite[2][29][77] = 1;dino_sprite[2][29][78] = 1;dino_sprite[2][29][79] = 1;dino_sprite[2][29][80] = 1;dino_sprite[2][29][81] = 1;dino_sprite[2][29][82] = 1;dino_sprite[2][29][83] = 1;dino_sprite[2][29][84] = 1;dino_sprite[2][29][85] = 1;dino_sprite[2][29][86] = 1;dino_sprite[2][29][87] = 1;dino_sprite[2][29][88] = 1;dino_sprite[2][29][89] = 1;dino_sprite[2][29][90] = 1;dino_sprite[2][29][91] = 1;dino_sprite[2][29][92] = 1;dino_sprite[2][29][93] = 1;dino_sprite[2][29][94] = 1;dino_sprite[2][29][95] = 1;dino_sprite[2][29][96] = 1;dino_sprite[2][29][97] = 1;dino_sprite[2][29][98] = 1;dino_sprite[2][29][99] = 1;dino_sprite[2][30][49] = 1;dino_sprite[2][30][50] = 1;dino_sprite[2][30][51] = 1;dino_sprite[2][30][52] = 1;dino_sprite[2][30][53] = 1;dino_sprite[2][30][54] = 1;dino_sprite[2][30][55] = 1;dino_sprite[2][30][56] = 1;dino_sprite[2][30][57] = 1;dino_sprite[2][30][58] = 1;dino_sprite[2][30][59] = 1;dino_sprite[2][30][60] = 1;dino_sprite[2][30][61] = 1;dino_sprite[2][30][62] = 1;dino_sprite[2][30][63] = 1;dino_sprite[2][30][64] = 1;dino_sprite[2][30][65] = 1;dino_sprite[2][30][66] = 1;dino_sprite[2][30][67] = 1;dino_sprite[2][30][68] = 1;dino_sprite[2][30][69] = 1;dino_sprite[2][30][70] = 1;dino_sprite[2][30][71] = 1;dino_sprite[2][30][72] = 1;dino_sprite[2][30][73] = 1;dino_sprite[2][30][74] = 1;dino_sprite[2][30][75] = 1;dino_sprite[2][30][76] = 1;dino_sprite[2][30][77] = 1;dino_sprite[2][30][78] = 1;dino_sprite[2][30][79] = 1;dino_sprite[2][30][80] = 1;dino_sprite[2][30][81] = 1;dino_sprite[2][30][82] = 1;dino_sprite[2][30][83] = 1;dino_sprite[2][30][84] = 1;dino_sprite[2][30][85] = 1;dino_sprite[2][30][86] = 1;dino_sprite[2][30][87] = 1;dino_sprite[2][30][88] = 1;dino_sprite[2][30][89] = 1;dino_sprite[2][30][90] = 1;dino_sprite[2][30][91] = 1;dino_sprite[2][30][92] = 1;dino_sprite[2][30][93] = 1;dino_sprite[2][30][94] = 1;dino_sprite[2][30][95] = 1;dino_sprite[2][30][96] = 1;dino_sprite[2][30][97] = 1;dino_sprite[2][30][98] = 1;dino_sprite[2][30][99] = 1;dino_sprite[2][31][44] = 1;dino_sprite[2][31][45] = 1;dino_sprite[2][31][46] = 1;dino_sprite[2][31][47] = 1;dino_sprite[2][31][48] = 1;dino_sprite[2][31][49] = 1;dino_sprite[2][31][50] = 1;dino_sprite[2][31][51] = 1;dino_sprite[2][31][52] = 1;dino_sprite[2][31][53] = 1;dino_sprite[2][31][54] = 1;dino_sprite[2][31][55] = 1;dino_sprite[2][31][56] = 1;dino_sprite[2][31][57] = 1;dino_sprite[2][31][58] = 1;dino_sprite[2][31][59] = 1;dino_sprite[2][31][60] = 1;dino_sprite[2][31][61] = 1;dino_sprite[2][31][62] = 1;dino_sprite[2][31][63] = 1;dino_sprite[2][31][64] = 1;dino_sprite[2][31][65] = 1;dino_sprite[2][31][66] = 1;dino_sprite[2][31][67] = 1;dino_sprite[2][31][68] = 1;dino_sprite[2][31][69] = 1;dino_sprite[2][31][70] = 1;dino_sprite[2][31][71] = 1;dino_sprite[2][31][72] = 1;dino_sprite[2][31][73] = 1;dino_sprite[2][31][74] = 1;dino_sprite[2][31][75] = 1;dino_sprite[2][31][76] = 1;dino_sprite[2][31][77] = 1;dino_sprite[2][31][78] = 1;dino_sprite[2][31][79] = 1;dino_sprite[2][31][80] = 1;dino_sprite[2][31][81] = 1;dino_sprite[2][31][82] = 1;dino_sprite[2][31][83] = 1;dino_sprite[2][31][84] = 1;dino_sprite[2][31][85] = 1;dino_sprite[2][31][86] = 1;dino_sprite[2][31][87] = 1;dino_sprite[2][31][88] = 1;dino_sprite[2][31][89] = 1;dino_sprite[2][31][90] = 1;dino_sprite[2][31][91] = 1;dino_sprite[2][31][92] = 1;dino_sprite[2][31][93] = 1;dino_sprite[2][31][94] = 1;dino_sprite[2][31][95] = 1;dino_sprite[2][31][96] = 1;dino_sprite[2][31][97] = 1;dino_sprite[2][31][98] = 1;dino_sprite[2][31][99] = 1;dino_sprite[2][32][44] = 1;dino_sprite[2][32][45] = 1;dino_sprite[2][32][46] = 1;dino_sprite[2][32][47] = 1;dino_sprite[2][32][48] = 1;dino_sprite[2][32][49] = 1;dino_sprite[2][32][50] = 1;dino_sprite[2][32][51] = 1;dino_sprite[2][32][52] = 1;dino_sprite[2][32][53] = 1;dino_sprite[2][32][54] = 1;dino_sprite[2][32][55] = 1;dino_sprite[2][32][56] = 1;dino_sprite[2][32][57] = 1;dino_sprite[2][32][58] = 1;dino_sprite[2][32][59] = 1;dino_sprite[2][32][60] = 1;dino_sprite[2][32][61] = 1;dino_sprite[2][32][62] = 1;dino_sprite[2][32][63] = 1;dino_sprite[2][32][64] = 1;dino_sprite[2][32][65] = 1;dino_sprite[2][32][66] = 1;dino_sprite[2][32][67] = 1;dino_sprite[2][32][68] = 1;dino_sprite[2][32][69] = 1;dino_sprite[2][32][70] = 1;dino_sprite[2][32][71] = 1;dino_sprite[2][32][72] = 1;dino_sprite[2][32][73] = 1;dino_sprite[2][32][74] = 1;dino_sprite[2][32][75] = 1;dino_sprite[2][32][76] = 1;dino_sprite[2][32][77] = 1;dino_sprite[2][32][78] = 1;dino_sprite[2][32][79] = 1;dino_sprite[2][32][80] = 1;dino_sprite[2][32][81] = 1;dino_sprite[2][32][82] = 1;dino_sprite[2][32][83] = 1;dino_sprite[2][32][84] = 1;dino_sprite[2][32][85] = 1;dino_sprite[2][32][86] = 1;dino_sprite[2][32][95] = 1;dino_sprite[2][32][96] = 1;dino_sprite[2][32][97] = 1;dino_sprite[2][32][98] = 1;dino_sprite[2][32][99] = 1;dino_sprite[2][33][44] = 1;dino_sprite[2][33][45] = 1;dino_sprite[2][33][46] = 1;dino_sprite[2][33][47] = 1;dino_sprite[2][33][48] = 1;dino_sprite[2][33][49] = 1;dino_sprite[2][33][50] = 1;dino_sprite[2][33][51] = 1;dino_sprite[2][33][52] = 1;dino_sprite[2][33][53] = 1;dino_sprite[2][33][54] = 1;dino_sprite[2][33][55] = 1;dino_sprite[2][33][56] = 1;dino_sprite[2][33][57] = 1;dino_sprite[2][33][58] = 1;dino_sprite[2][33][59] = 1;dino_sprite[2][33][60] = 1;dino_sprite[2][33][61] = 1;dino_sprite[2][33][62] = 1;dino_sprite[2][33][63] = 1;dino_sprite[2][33][64] = 1;dino_sprite[2][33][65] = 1;dino_sprite[2][33][66] = 1;dino_sprite[2][33][67] = 1;dino_sprite[2][33][68] = 1;dino_sprite[2][33][69] = 1;dino_sprite[2][33][70] = 1;dino_sprite[2][33][71] = 1;dino_sprite[2][33][72] = 1;dino_sprite[2][33][73] = 1;dino_sprite[2][33][74] = 1;dino_sprite[2][33][75] = 1;dino_sprite[2][33][76] = 1;dino_sprite[2][33][77] = 1;dino_sprite[2][33][78] = 1;dino_sprite[2][33][79] = 1;dino_sprite[2][33][80] = 1;dino_sprite[2][33][81] = 1;dino_sprite[2][33][82] = 1;dino_sprite[2][33][83] = 1;dino_sprite[2][33][84] = 1;dino_sprite[2][33][85] = 1;dino_sprite[2][33][86] = 1;dino_sprite[2][33][95] = 1;dino_sprite[2][33][96] = 1;dino_sprite[2][33][97] = 1;dino_sprite[2][33][98] = 1;dino_sprite[2][33][99] = 1;dino_sprite[2][34][44] = 1;dino_sprite[2][34][45] = 1;dino_sprite[2][34][46] = 1;dino_sprite[2][34][47] = 1;dino_sprite[2][34][48] = 1;dino_sprite[2][34][49] = 1;dino_sprite[2][34][50] = 1;dino_sprite[2][34][51] = 1;dino_sprite[2][34][52] = 1;dino_sprite[2][34][53] = 1;dino_sprite[2][34][54] = 1;dino_sprite[2][34][55] = 1;dino_sprite[2][34][56] = 1;dino_sprite[2][34][57] = 1;dino_sprite[2][34][58] = 1;dino_sprite[2][34][59] = 1;dino_sprite[2][34][60] = 1;dino_sprite[2][34][61] = 1;dino_sprite[2][34][62] = 1;dino_sprite[2][34][63] = 1;dino_sprite[2][34][64] = 1;dino_sprite[2][34][65] = 1;dino_sprite[2][34][66] = 1;dino_sprite[2][34][67] = 1;dino_sprite[2][34][68] = 1;dino_sprite[2][34][69] = 1;dino_sprite[2][34][70] = 1;dino_sprite[2][34][71] = 1;dino_sprite[2][34][72] = 1;dino_sprite[2][34][73] = 1;dino_sprite[2][34][74] = 1;dino_sprite[2][34][75] = 1;dino_sprite[2][34][76] = 1;dino_sprite[2][34][77] = 1;dino_sprite[2][34][78] = 1;dino_sprite[2][34][79] = 1;dino_sprite[2][34][80] = 1;dino_sprite[2][34][81] = 1;dino_sprite[2][34][82] = 1;dino_sprite[2][34][83] = 1;dino_sprite[2][34][84] = 1;dino_sprite[2][34][85] = 1;dino_sprite[2][34][86] = 1;dino_sprite[2][34][95] = 1;dino_sprite[2][34][96] = 1;dino_sprite[2][34][97] = 1;dino_sprite[2][34][98] = 1;dino_sprite[2][34][99] = 1;dino_sprite[2][35][44] = 1;dino_sprite[2][35][45] = 1;dino_sprite[2][35][46] = 1;dino_sprite[2][35][47] = 1;dino_sprite[2][35][48] = 1;dino_sprite[2][35][49] = 1;dino_sprite[2][35][50] = 1;dino_sprite[2][35][51] = 1;dino_sprite[2][35][52] = 1;dino_sprite[2][35][53] = 1;dino_sprite[2][35][54] = 1;dino_sprite[2][35][55] = 1;dino_sprite[2][35][56] = 1;dino_sprite[2][35][57] = 1;dino_sprite[2][35][58] = 1;dino_sprite[2][35][59] = 1;dino_sprite[2][35][60] = 1;dino_sprite[2][35][61] = 1;dino_sprite[2][35][62] = 1;dino_sprite[2][35][63] = 1;dino_sprite[2][35][64] = 1;dino_sprite[2][35][65] = 1;dino_sprite[2][35][66] = 1;dino_sprite[2][35][67] = 1;dino_sprite[2][35][68] = 1;dino_sprite[2][35][69] = 1;dino_sprite[2][35][70] = 1;dino_sprite[2][35][71] = 1;dino_sprite[2][35][72] = 1;dino_sprite[2][35][73] = 1;dino_sprite[2][35][74] = 1;dino_sprite[2][35][75] = 1;dino_sprite[2][35][76] = 1;dino_sprite[2][35][77] = 1;dino_sprite[2][35][78] = 1;dino_sprite[2][35][79] = 1;dino_sprite[2][35][80] = 1;dino_sprite[2][35][81] = 1;dino_sprite[2][35][82] = 1;dino_sprite[2][35][83] = 1;dino_sprite[2][35][84] = 1;dino_sprite[2][35][85] = 1;dino_sprite[2][35][86] = 1;dino_sprite[2][35][95] = 1;dino_sprite[2][35][96] = 1;dino_sprite[2][35][97] = 1;dino_sprite[2][35][98] = 1;dino_sprite[2][35][99] = 1;dino_sprite[2][36][44] = 1;dino_sprite[2][36][45] = 1;dino_sprite[2][36][46] = 1;dino_sprite[2][36][47] = 1;dino_sprite[2][36][48] = 1;dino_sprite[2][36][49] = 1;dino_sprite[2][36][50] = 1;dino_sprite[2][36][51] = 1;dino_sprite[2][36][52] = 1;dino_sprite[2][36][53] = 1;dino_sprite[2][36][54] = 1;dino_sprite[2][36][55] = 1;dino_sprite[2][36][56] = 1;dino_sprite[2][36][57] = 1;dino_sprite[2][36][58] = 1;dino_sprite[2][36][59] = 1;dino_sprite[2][36][60] = 1;dino_sprite[2][36][61] = 1;dino_sprite[2][36][62] = 1;dino_sprite[2][36][63] = 1;dino_sprite[2][36][64] = 1;dino_sprite[2][36][65] = 1;dino_sprite[2][36][66] = 1;dino_sprite[2][36][67] = 1;dino_sprite[2][36][68] = 1;dino_sprite[2][36][69] = 1;dino_sprite[2][36][70] = 1;dino_sprite[2][36][71] = 1;dino_sprite[2][36][72] = 1;dino_sprite[2][36][73] = 1;dino_sprite[2][36][74] = 1;dino_sprite[2][36][75] = 1;dino_sprite[2][36][76] = 1;dino_sprite[2][36][77] = 1;dino_sprite[2][36][78] = 1;dino_sprite[2][36][79] = 1;dino_sprite[2][36][80] = 1;dino_sprite[2][36][81] = 1;dino_sprite[2][36][82] = 1;dino_sprite[2][36][83] = 1;dino_sprite[2][36][84] = 1;dino_sprite[2][36][85] = 1;dino_sprite[2][36][86] = 1;dino_sprite[2][36][95] = 1;dino_sprite[2][36][96] = 1;dino_sprite[2][36][97] = 1;dino_sprite[2][36][98] = 1;dino_sprite[2][36][99] = 1;dino_sprite[2][37][44] = 1;dino_sprite[2][37][45] = 1;dino_sprite[2][37][46] = 1;dino_sprite[2][37][47] = 1;dino_sprite[2][37][48] = 1;dino_sprite[2][37][49] = 1;dino_sprite[2][37][50] = 1;dino_sprite[2][37][51] = 1;dino_sprite[2][37][52] = 1;dino_sprite[2][37][53] = 1;dino_sprite[2][37][54] = 1;dino_sprite[2][37][55] = 1;dino_sprite[2][37][56] = 1;dino_sprite[2][37][57] = 1;dino_sprite[2][37][58] = 1;dino_sprite[2][37][59] = 1;dino_sprite[2][37][60] = 1;dino_sprite[2][37][61] = 1;dino_sprite[2][37][62] = 1;dino_sprite[2][37][63] = 1;dino_sprite[2][37][64] = 1;dino_sprite[2][37][65] = 1;dino_sprite[2][37][66] = 1;dino_sprite[2][37][67] = 1;dino_sprite[2][37][68] = 1;dino_sprite[2][37][69] = 1;dino_sprite[2][37][70] = 1;dino_sprite[2][37][71] = 1;dino_sprite[2][37][72] = 1;dino_sprite[2][37][73] = 1;dino_sprite[2][37][74] = 1;dino_sprite[2][37][75] = 1;dino_sprite[2][37][76] = 1;dino_sprite[2][37][77] = 1;dino_sprite[2][37][78] = 1;dino_sprite[2][37][79] = 1;dino_sprite[2][37][80] = 1;dino_sprite[2][37][81] = 1;dino_sprite[2][37][82] = 1;dino_sprite[2][37][83] = 1;dino_sprite[2][37][84] = 1;dino_sprite[2][37][85] = 1;dino_sprite[2][37][86] = 1;dino_sprite[2][38][44] = 1;dino_sprite[2][38][45] = 1;dino_sprite[2][38][46] = 1;dino_sprite[2][38][47] = 1;dino_sprite[2][38][48] = 1;dino_sprite[2][38][49] = 1;dino_sprite[2][38][50] = 1;dino_sprite[2][38][51] = 1;dino_sprite[2][38][52] = 1;dino_sprite[2][38][53] = 1;dino_sprite[2][38][54] = 1;dino_sprite[2][38][55] = 1;dino_sprite[2][38][56] = 1;dino_sprite[2][38][57] = 1;dino_sprite[2][38][58] = 1;dino_sprite[2][38][59] = 1;dino_sprite[2][38][60] = 1;dino_sprite[2][38][61] = 1;dino_sprite[2][38][62] = 1;dino_sprite[2][38][63] = 1;dino_sprite[2][38][64] = 1;dino_sprite[2][38][65] = 1;dino_sprite[2][38][66] = 1;dino_sprite[2][38][67] = 1;dino_sprite[2][38][68] = 1;dino_sprite[2][38][69] = 1;dino_sprite[2][38][70] = 1;dino_sprite[2][38][71] = 1;dino_sprite[2][38][72] = 1;dino_sprite[2][38][73] = 1;dino_sprite[2][38][74] = 1;dino_sprite[2][38][75] = 1;dino_sprite[2][38][76] = 1;dino_sprite[2][38][77] = 1;dino_sprite[2][38][78] = 1;dino_sprite[2][38][79] = 1;dino_sprite[2][38][80] = 1;dino_sprite[2][38][81] = 1;dino_sprite[2][38][82] = 1;dino_sprite[2][38][83] = 1;dino_sprite[2][38][84] = 1;dino_sprite[2][38][85] = 1;dino_sprite[2][38][86] = 1;dino_sprite[2][39][39] = 1;dino_sprite[2][39][40] = 1;dino_sprite[2][39][41] = 1;dino_sprite[2][39][42] = 1;dino_sprite[2][39][43] = 1;dino_sprite[2][39][44] = 1;dino_sprite[2][39][45] = 1;dino_sprite[2][39][46] = 1;dino_sprite[2][39][47] = 1;dino_sprite[2][39][48] = 1;dino_sprite[2][39][49] = 1;dino_sprite[2][39][50] = 1;dino_sprite[2][39][51] = 1;dino_sprite[2][39][52] = 1;dino_sprite[2][39][53] = 1;dino_sprite[2][39][54] = 1;dino_sprite[2][39][55] = 1;dino_sprite[2][39][56] = 1;dino_sprite[2][39][57] = 1;dino_sprite[2][39][58] = 1;dino_sprite[2][39][59] = 1;dino_sprite[2][39][60] = 1;dino_sprite[2][39][61] = 1;dino_sprite[2][39][62] = 1;dino_sprite[2][39][63] = 1;dino_sprite[2][39][64] = 1;dino_sprite[2][39][65] = 1;dino_sprite[2][39][66] = 1;dino_sprite[2][39][67] = 1;dino_sprite[2][39][68] = 1;dino_sprite[2][39][69] = 1;dino_sprite[2][39][70] = 1;dino_sprite[2][39][71] = 1;dino_sprite[2][39][72] = 1;dino_sprite[2][39][73] = 1;dino_sprite[2][39][74] = 1;dino_sprite[2][39][75] = 1;dino_sprite[2][39][76] = 1;dino_sprite[2][39][77] = 1;dino_sprite[2][39][78] = 1;dino_sprite[2][39][79] = 1;dino_sprite[2][39][80] = 1;dino_sprite[2][39][81] = 1;dino_sprite[2][39][82] = 1;dino_sprite[2][39][83] = 1;dino_sprite[2][39][84] = 1;dino_sprite[2][39][85] = 1;dino_sprite[2][39][86] = 1;dino_sprite[2][40][39] = 1;dino_sprite[2][40][40] = 1;dino_sprite[2][40][41] = 1;dino_sprite[2][40][42] = 1;dino_sprite[2][40][43] = 1;dino_sprite[2][40][44] = 1;dino_sprite[2][40][45] = 1;dino_sprite[2][40][46] = 1;dino_sprite[2][40][47] = 1;dino_sprite[2][40][48] = 1;dino_sprite[2][40][49] = 1;dino_sprite[2][40][50] = 1;dino_sprite[2][40][51] = 1;dino_sprite[2][40][52] = 1;dino_sprite[2][40][53] = 1;dino_sprite[2][40][54] = 1;dino_sprite[2][40][55] = 1;dino_sprite[2][40][56] = 1;dino_sprite[2][40][57] = 1;dino_sprite[2][40][58] = 1;dino_sprite[2][40][59] = 1;dino_sprite[2][40][60] = 1;dino_sprite[2][40][61] = 1;dino_sprite[2][40][62] = 1;dino_sprite[2][40][63] = 1;dino_sprite[2][40][64] = 1;dino_sprite[2][40][65] = 1;dino_sprite[2][40][66] = 1;dino_sprite[2][40][67] = 1;dino_sprite[2][40][68] = 1;dino_sprite[2][40][69] = 1;dino_sprite[2][40][70] = 1;dino_sprite[2][40][71] = 1;dino_sprite[2][40][72] = 1;dino_sprite[2][40][73] = 1;dino_sprite[2][40][74] = 1;dino_sprite[2][40][75] = 1;dino_sprite[2][40][76] = 1;dino_sprite[2][40][77] = 1;dino_sprite[2][40][78] = 1;dino_sprite[2][40][79] = 1;dino_sprite[2][40][80] = 1;dino_sprite[2][40][81] = 1;dino_sprite[2][40][82] = 1;dino_sprite[2][40][83] = 1;dino_sprite[2][40][84] = 1;dino_sprite[2][40][85] = 1;dino_sprite[2][40][86] = 1;dino_sprite[2][41][39] = 1;dino_sprite[2][41][40] = 1;dino_sprite[2][41][41] = 1;dino_sprite[2][41][42] = 1;dino_sprite[2][41][43] = 1;dino_sprite[2][41][44] = 1;dino_sprite[2][41][45] = 1;dino_sprite[2][41][46] = 1;dino_sprite[2][41][47] = 1;dino_sprite[2][41][48] = 1;dino_sprite[2][41][49] = 1;dino_sprite[2][41][50] = 1;dino_sprite[2][41][51] = 1;dino_sprite[2][41][52] = 1;dino_sprite[2][41][53] = 1;dino_sprite[2][41][54] = 1;dino_sprite[2][41][55] = 1;dino_sprite[2][41][56] = 1;dino_sprite[2][41][57] = 1;dino_sprite[2][41][58] = 1;dino_sprite[2][41][59] = 1;dino_sprite[2][41][60] = 1;dino_sprite[2][41][61] = 1;dino_sprite[2][41][62] = 1;dino_sprite[2][41][63] = 1;dino_sprite[2][41][64] = 1;dino_sprite[2][41][65] = 1;dino_sprite[2][41][66] = 1;dino_sprite[2][41][67] = 1;dino_sprite[2][41][68] = 1;dino_sprite[2][41][69] = 1;dino_sprite[2][41][70] = 1;dino_sprite[2][41][71] = 1;dino_sprite[2][41][72] = 1;dino_sprite[2][41][73] = 1;dino_sprite[2][41][74] = 1;dino_sprite[2][41][75] = 1;dino_sprite[2][41][76] = 1;dino_sprite[2][41][77] = 1;dino_sprite[2][41][78] = 1;dino_sprite[2][41][79] = 1;dino_sprite[2][41][80] = 1;dino_sprite[2][41][81] = 1;dino_sprite[2][41][82] = 1;dino_sprite[2][42][39] = 1;dino_sprite[2][42][40] = 1;dino_sprite[2][42][41] = 1;dino_sprite[2][42][42] = 1;dino_sprite[2][42][43] = 1;dino_sprite[2][42][44] = 1;dino_sprite[2][42][45] = 1;dino_sprite[2][42][46] = 1;dino_sprite[2][42][47] = 1;dino_sprite[2][42][48] = 1;dino_sprite[2][42][49] = 1;dino_sprite[2][42][50] = 1;dino_sprite[2][42][51] = 1;dino_sprite[2][42][52] = 1;dino_sprite[2][42][53] = 1;dino_sprite[2][42][54] = 1;dino_sprite[2][42][55] = 1;dino_sprite[2][42][56] = 1;dino_sprite[2][42][57] = 1;dino_sprite[2][42][58] = 1;dino_sprite[2][42][59] = 1;dino_sprite[2][42][60] = 1;dino_sprite[2][42][61] = 1;dino_sprite[2][42][62] = 1;dino_sprite[2][42][63] = 1;dino_sprite[2][42][64] = 1;dino_sprite[2][42][65] = 1;dino_sprite[2][42][66] = 1;dino_sprite[2][42][67] = 1;dino_sprite[2][42][68] = 1;dino_sprite[2][42][69] = 1;dino_sprite[2][42][70] = 1;dino_sprite[2][42][71] = 1;dino_sprite[2][42][72] = 1;dino_sprite[2][42][73] = 1;dino_sprite[2][42][74] = 1;dino_sprite[2][42][75] = 1;dino_sprite[2][42][76] = 1;dino_sprite[2][42][77] = 1;dino_sprite[2][42][78] = 1;dino_sprite[2][42][79] = 1;dino_sprite[2][42][80] = 1;dino_sprite[2][42][81] = 1;dino_sprite[2][42][82] = 1;dino_sprite[2][43][39] = 1;dino_sprite[2][43][40] = 1;dino_sprite[2][43][41] = 1;dino_sprite[2][43][42] = 1;dino_sprite[2][43][43] = 1;dino_sprite[2][43][44] = 1;dino_sprite[2][43][45] = 1;dino_sprite[2][43][46] = 1;dino_sprite[2][43][47] = 1;dino_sprite[2][43][48] = 1;dino_sprite[2][43][49] = 1;dino_sprite[2][43][50] = 1;dino_sprite[2][43][51] = 1;dino_sprite[2][43][52] = 1;dino_sprite[2][43][53] = 1;dino_sprite[2][43][54] = 1;dino_sprite[2][43][55] = 1;dino_sprite[2][43][56] = 1;dino_sprite[2][43][57] = 1;dino_sprite[2][43][58] = 1;dino_sprite[2][43][59] = 1;dino_sprite[2][43][60] = 1;dino_sprite[2][43][61] = 1;dino_sprite[2][43][62] = 1;dino_sprite[2][43][63] = 1;dino_sprite[2][43][64] = 1;dino_sprite[2][43][65] = 1;dino_sprite[2][43][66] = 1;dino_sprite[2][43][67] = 1;dino_sprite[2][43][68] = 1;dino_sprite[2][43][69] = 1;dino_sprite[2][43][70] = 1;dino_sprite[2][43][71] = 1;dino_sprite[2][43][72] = 1;dino_sprite[2][43][73] = 1;dino_sprite[2][43][74] = 1;dino_sprite[2][43][75] = 1;dino_sprite[2][43][76] = 1;dino_sprite[2][43][77] = 1;dino_sprite[2][43][78] = 1;dino_sprite[2][43][79] = 1;dino_sprite[2][43][80] = 1;dino_sprite[2][43][81] = 1;dino_sprite[2][43][82] = 1;dino_sprite[2][44][39] = 1;dino_sprite[2][44][40] = 1;dino_sprite[2][44][41] = 1;dino_sprite[2][44][42] = 1;dino_sprite[2][44][43] = 1;dino_sprite[2][44][44] = 1;dino_sprite[2][44][45] = 1;dino_sprite[2][44][46] = 1;dino_sprite[2][44][47] = 1;dino_sprite[2][44][48] = 1;dino_sprite[2][44][49] = 1;dino_sprite[2][44][50] = 1;dino_sprite[2][44][51] = 1;dino_sprite[2][44][52] = 1;dino_sprite[2][44][53] = 1;dino_sprite[2][44][54] = 1;dino_sprite[2][44][55] = 1;dino_sprite[2][44][56] = 1;dino_sprite[2][44][57] = 1;dino_sprite[2][44][58] = 1;dino_sprite[2][44][59] = 1;dino_sprite[2][44][60] = 1;dino_sprite[2][44][61] = 1;dino_sprite[2][44][62] = 1;dino_sprite[2][44][63] = 1;dino_sprite[2][44][64] = 1;dino_sprite[2][44][65] = 1;dino_sprite[2][44][66] = 1;dino_sprite[2][44][67] = 1;dino_sprite[2][44][68] = 1;dino_sprite[2][44][69] = 1;dino_sprite[2][44][70] = 1;dino_sprite[2][44][71] = 1;dino_sprite[2][44][72] = 1;dino_sprite[2][44][73] = 1;dino_sprite[2][44][74] = 1;dino_sprite[2][44][75] = 1;dino_sprite[2][44][76] = 1;dino_sprite[2][44][77] = 1;dino_sprite[2][44][78] = 1;dino_sprite[2][44][79] = 1;dino_sprite[2][44][80] = 1;dino_sprite[2][44][81] = 1;dino_sprite[2][44][82] = 1;dino_sprite[2][45][35] = 1;dino_sprite[2][45][36] = 1;dino_sprite[2][45][37] = 1;dino_sprite[2][45][39] = 1;dino_sprite[2][45][40] = 1;dino_sprite[2][45][41] = 1;dino_sprite[2][45][42] = 1;dino_sprite[2][45][43] = 1;dino_sprite[2][45][44] = 1;dino_sprite[2][45][45] = 1;dino_sprite[2][45][46] = 1;dino_sprite[2][45][47] = 1;dino_sprite[2][45][48] = 1;dino_sprite[2][45][49] = 1;dino_sprite[2][45][50] = 1;dino_sprite[2][45][51] = 1;dino_sprite[2][45][52] = 1;dino_sprite[2][45][53] = 1;dino_sprite[2][45][54] = 1;dino_sprite[2][45][55] = 1;dino_sprite[2][45][56] = 1;dino_sprite[2][45][57] = 1;dino_sprite[2][45][58] = 1;dino_sprite[2][45][59] = 1;dino_sprite[2][45][60] = 1;dino_sprite[2][45][61] = 1;dino_sprite[2][45][62] = 1;dino_sprite[2][45][63] = 1;dino_sprite[2][45][64] = 1;dino_sprite[2][45][65] = 1;dino_sprite[2][45][66] = 1;dino_sprite[2][45][67] = 1;dino_sprite[2][45][68] = 1;dino_sprite[2][45][69] = 1;dino_sprite[2][45][70] = 1;dino_sprite[2][45][71] = 1;dino_sprite[2][45][72] = 1;dino_sprite[2][45][73] = 1;dino_sprite[2][45][74] = 1;dino_sprite[2][45][75] = 1;dino_sprite[2][45][76] = 1;dino_sprite[2][45][77] = 1;dino_sprite[2][45][78] = 1;dino_sprite[2][45][79] = 1;dino_sprite[2][45][80] = 1;dino_sprite[2][45][81] = 1;dino_sprite[2][45][82] = 1;dino_sprite[2][45][84] = 1;dino_sprite[2][45][85] = 1;dino_sprite[2][45][86] = 1;dino_sprite[2][46][35] = 1;dino_sprite[2][46][36] = 1;dino_sprite[2][46][37] = 1;dino_sprite[2][46][38] = 1;dino_sprite[2][46][39] = 1;dino_sprite[2][46][40] = 1;dino_sprite[2][46][41] = 1;dino_sprite[2][46][42] = 1;dino_sprite[2][46][43] = 1;dino_sprite[2][46][44] = 1;dino_sprite[2][46][45] = 1;dino_sprite[2][46][46] = 1;dino_sprite[2][46][47] = 1;dino_sprite[2][46][48] = 1;dino_sprite[2][46][49] = 1;dino_sprite[2][46][50] = 1;dino_sprite[2][46][51] = 1;dino_sprite[2][46][52] = 1;dino_sprite[2][46][53] = 1;dino_sprite[2][46][54] = 1;dino_sprite[2][46][55] = 1;dino_sprite[2][46][56] = 1;dino_sprite[2][46][57] = 1;dino_sprite[2][46][58] = 1;dino_sprite[2][46][59] = 1;dino_sprite[2][46][60] = 1;dino_sprite[2][46][61] = 1;dino_sprite[2][46][62] = 1;dino_sprite[2][46][63] = 1;dino_sprite[2][46][64] = 1;dino_sprite[2][46][65] = 1;dino_sprite[2][46][66] = 1;dino_sprite[2][46][67] = 1;dino_sprite[2][46][68] = 1;dino_sprite[2][46][69] = 1;dino_sprite[2][46][70] = 1;dino_sprite[2][46][71] = 1;dino_sprite[2][46][72] = 1;dino_sprite[2][46][73] = 1;dino_sprite[2][46][74] = 1;dino_sprite[2][46][75] = 1;dino_sprite[2][46][76] = 1;dino_sprite[2][46][77] = 1;dino_sprite[2][46][78] = 1;dino_sprite[2][46][79] = 1;dino_sprite[2][46][80] = 1;dino_sprite[2][46][81] = 1;dino_sprite[2][46][82] = 1;dino_sprite[2][46][83] = 1;dino_sprite[2][46][84] = 1;dino_sprite[2][46][85] = 1;dino_sprite[2][46][86] = 1;dino_sprite[2][47][35] = 1;dino_sprite[2][47][36] = 1;dino_sprite[2][47][37] = 1;dino_sprite[2][47][38] = 1;dino_sprite[2][47][39] = 1;dino_sprite[2][47][40] = 1;dino_sprite[2][47][41] = 1;dino_sprite[2][47][42] = 1;dino_sprite[2][47][43] = 1;dino_sprite[2][47][44] = 1;dino_sprite[2][47][45] = 1;dino_sprite[2][47][46] = 1;dino_sprite[2][47][47] = 1;dino_sprite[2][47][48] = 1;dino_sprite[2][47][49] = 1;dino_sprite[2][47][50] = 1;dino_sprite[2][47][51] = 1;dino_sprite[2][47][52] = 1;dino_sprite[2][47][53] = 1;dino_sprite[2][47][54] = 1;dino_sprite[2][47][55] = 1;dino_sprite[2][47][56] = 1;dino_sprite[2][47][57] = 1;dino_sprite[2][47][58] = 1;dino_sprite[2][47][59] = 1;dino_sprite[2][47][60] = 1;dino_sprite[2][47][61] = 1;dino_sprite[2][47][62] = 1;dino_sprite[2][47][63] = 1;dino_sprite[2][47][64] = 1;dino_sprite[2][47][65] = 1;dino_sprite[2][47][66] = 1;dino_sprite[2][47][67] = 1;dino_sprite[2][47][68] = 1;dino_sprite[2][47][69] = 1;dino_sprite[2][47][70] = 1;dino_sprite[2][47][71] = 1;dino_sprite[2][47][72] = 1;dino_sprite[2][47][73] = 1;dino_sprite[2][47][74] = 1;dino_sprite[2][47][75] = 1;dino_sprite[2][47][76] = 1;dino_sprite[2][47][77] = 1;dino_sprite[2][47][78] = 1;dino_sprite[2][47][79] = 1;dino_sprite[2][47][80] = 1;dino_sprite[2][47][81] = 1;dino_sprite[2][47][82] = 1;dino_sprite[2][47][83] = 1;dino_sprite[2][47][84] = 1;dino_sprite[2][47][85] = 1;dino_sprite[2][47][86] = 1;dino_sprite[2][48][35] = 1;dino_sprite[2][48][36] = 1;dino_sprite[2][48][37] = 1;dino_sprite[2][48][38] = 1;dino_sprite[2][48][39] = 1;dino_sprite[2][48][40] = 1;dino_sprite[2][48][41] = 1;dino_sprite[2][48][42] = 1;dino_sprite[2][48][43] = 1;dino_sprite[2][48][44] = 1;dino_sprite[2][48][45] = 1;dino_sprite[2][48][46] = 1;dino_sprite[2][48][47] = 1;dino_sprite[2][48][48] = 1;dino_sprite[2][48][49] = 1;dino_sprite[2][48][50] = 1;dino_sprite[2][48][51] = 1;dino_sprite[2][48][52] = 1;dino_sprite[2][48][53] = 1;dino_sprite[2][48][54] = 1;dino_sprite[2][48][55] = 1;dino_sprite[2][48][56] = 1;dino_sprite[2][48][57] = 1;dino_sprite[2][48][58] = 1;dino_sprite[2][48][59] = 1;dino_sprite[2][48][60] = 1;dino_sprite[2][48][61] = 1;dino_sprite[2][48][62] = 1;dino_sprite[2][48][63] = 1;dino_sprite[2][48][64] = 1;dino_sprite[2][48][65] = 1;dino_sprite[2][48][66] = 1;dino_sprite[2][48][67] = 1;dino_sprite[2][48][68] = 1;dino_sprite[2][48][69] = 1;dino_sprite[2][48][70] = 1;dino_sprite[2][48][71] = 1;dino_sprite[2][48][72] = 1;dino_sprite[2][48][73] = 1;dino_sprite[2][48][74] = 1;dino_sprite[2][48][75] = 1;dino_sprite[2][48][76] = 1;dino_sprite[2][48][77] = 1;dino_sprite[2][48][78] = 1;dino_sprite[2][48][79] = 1;dino_sprite[2][48][80] = 1;dino_sprite[2][48][81] = 1;dino_sprite[2][48][82] = 1;dino_sprite[2][48][83] = 1;dino_sprite[2][48][84] = 1;dino_sprite[2][48][85] = 1;dino_sprite[2][48][86] = 1;dino_sprite[2][49][35] = 1;dino_sprite[2][49][36] = 1;dino_sprite[2][49][37] = 1;dino_sprite[2][49][38] = 1;dino_sprite[2][49][39] = 1;dino_sprite[2][49][40] = 1;dino_sprite[2][49][41] = 1;dino_sprite[2][49][42] = 1;dino_sprite[2][49][43] = 1;dino_sprite[2][49][44] = 1;dino_sprite[2][49][45] = 1;dino_sprite[2][49][46] = 1;dino_sprite[2][49][47] = 1;dino_sprite[2][49][48] = 1;dino_sprite[2][49][49] = 1;dino_sprite[2][49][50] = 1;dino_sprite[2][49][51] = 1;dino_sprite[2][49][52] = 1;dino_sprite[2][49][53] = 1;dino_sprite[2][49][54] = 1;dino_sprite[2][49][55] = 1;dino_sprite[2][49][56] = 1;dino_sprite[2][49][57] = 1;dino_sprite[2][49][58] = 1;dino_sprite[2][49][59] = 1;dino_sprite[2][49][60] = 1;dino_sprite[2][49][61] = 1;dino_sprite[2][49][62] = 1;dino_sprite[2][49][63] = 1;dino_sprite[2][49][64] = 1;dino_sprite[2][49][65] = 1;dino_sprite[2][49][66] = 1;dino_sprite[2][49][67] = 1;dino_sprite[2][49][68] = 1;dino_sprite[2][49][69] = 1;dino_sprite[2][49][70] = 1;dino_sprite[2][49][71] = 1;dino_sprite[2][49][72] = 1;dino_sprite[2][49][73] = 1;dino_sprite[2][49][74] = 1;dino_sprite[2][49][75] = 1;dino_sprite[2][49][76] = 1;dino_sprite[2][49][77] = 1;dino_sprite[2][49][78] = 1;dino_sprite[2][49][79] = 1;dino_sprite[2][49][80] = 1;dino_sprite[2][49][81] = 1;dino_sprite[2][49][82] = 1;dino_sprite[2][49][83] = 1;dino_sprite[2][49][84] = 1;dino_sprite[2][49][85] = 1;dino_sprite[2][49][86] = 1;dino_sprite[2][50][35] = 1;dino_sprite[2][50][36] = 1;dino_sprite[2][50][37] = 1;dino_sprite[2][50][38] = 1;dino_sprite[2][50][39] = 1;dino_sprite[2][50][40] = 1;dino_sprite[2][50][41] = 1;dino_sprite[2][50][42] = 1;dino_sprite[2][50][43] = 1;dino_sprite[2][50][44] = 1;dino_sprite[2][50][45] = 1;dino_sprite[2][50][46] = 1;dino_sprite[2][50][47] = 1;dino_sprite[2][50][48] = 1;dino_sprite[2][50][49] = 1;dino_sprite[2][50][50] = 1;dino_sprite[2][50][51] = 1;dino_sprite[2][50][52] = 1;dino_sprite[2][50][53] = 1;dino_sprite[2][50][54] = 1;dino_sprite[2][50][55] = 1;dino_sprite[2][50][56] = 1;dino_sprite[2][50][57] = 1;dino_sprite[2][50][58] = 1;dino_sprite[2][50][59] = 1;dino_sprite[2][50][60] = 1;dino_sprite[2][50][61] = 1;dino_sprite[2][50][62] = 1;dino_sprite[2][50][63] = 1;dino_sprite[2][50][64] = 1;dino_sprite[2][50][65] = 1;dino_sprite[2][50][66] = 1;dino_sprite[2][50][67] = 1;dino_sprite[2][50][68] = 1;dino_sprite[2][50][69] = 1;dino_sprite[2][50][70] = 1;dino_sprite[2][50][71] = 1;dino_sprite[2][50][72] = 1;dino_sprite[2][50][73] = 1;dino_sprite[2][50][74] = 1;dino_sprite[2][50][75] = 1;dino_sprite[2][50][76] = 1;dino_sprite[2][50][77] = 1;dino_sprite[2][50][78] = 1;dino_sprite[2][50][79] = 1;dino_sprite[2][50][80] = 1;dino_sprite[2][50][81] = 1;dino_sprite[2][50][82] = 1;dino_sprite[2][50][83] = 1;dino_sprite[2][50][84] = 1;dino_sprite[2][50][85] = 1;dino_sprite[2][50][86] = 1;dino_sprite[2][50][88] = 1;dino_sprite[2][50][89] = 1;dino_sprite[2][50][90] = 1;dino_sprite[2][50][91] = 1;dino_sprite[2][50][92] = 1;dino_sprite[2][51][3] = 1;dino_sprite[2][51][4] = 1;dino_sprite[2][51][5] = 1;dino_sprite[2][51][6] = 1;dino_sprite[2][51][7] = 1;dino_sprite[2][51][8] = 1;dino_sprite[2][51][9] = 1;dino_sprite[2][51][10] = 1;dino_sprite[2][51][11] = 1;dino_sprite[2][51][12] = 1;dino_sprite[2][51][13] = 1;dino_sprite[2][51][14] = 1;dino_sprite[2][51][15] = 1;dino_sprite[2][51][16] = 1;dino_sprite[2][51][17] = 1;dino_sprite[2][51][18] = 1;dino_sprite[2][51][19] = 1;dino_sprite[2][51][20] = 1;dino_sprite[2][51][21] = 1;dino_sprite[2][51][22] = 1;dino_sprite[2][51][23] = 1;dino_sprite[2][51][24] = 1;dino_sprite[2][51][25] = 1;dino_sprite[2][51][26] = 1;dino_sprite[2][51][27] = 1;dino_sprite[2][51][28] = 1;dino_sprite[2][51][29] = 1;dino_sprite[2][51][30] = 1;dino_sprite[2][51][31] = 1;dino_sprite[2][51][32] = 1;dino_sprite[2][51][33] = 1;dino_sprite[2][51][34] = 1;dino_sprite[2][51][35] = 1;dino_sprite[2][51][36] = 1;dino_sprite[2][51][37] = 1;dino_sprite[2][51][38] = 1;dino_sprite[2][51][39] = 1;dino_sprite[2][51][40] = 1;dino_sprite[2][51][41] = 1;dino_sprite[2][51][42] = 1;dino_sprite[2][51][43] = 1;dino_sprite[2][51][44] = 1;dino_sprite[2][51][45] = 1;dino_sprite[2][51][46] = 1;dino_sprite[2][51][47] = 1;dino_sprite[2][51][48] = 1;dino_sprite[2][51][49] = 1;dino_sprite[2][51][50] = 1;dino_sprite[2][51][51] = 1;dino_sprite[2][51][52] = 1;dino_sprite[2][51][53] = 1;dino_sprite[2][51][54] = 1;dino_sprite[2][51][55] = 1;dino_sprite[2][51][56] = 1;dino_sprite[2][51][57] = 1;dino_sprite[2][51][58] = 1;dino_sprite[2][51][59] = 1;dino_sprite[2][51][60] = 1;dino_sprite[2][51][61] = 1;dino_sprite[2][51][62] = 1;dino_sprite[2][51][63] = 1;dino_sprite[2][51][64] = 1;dino_sprite[2][51][65] = 1;dino_sprite[2][51][66] = 1;dino_sprite[2][51][67] = 1;dino_sprite[2][51][68] = 1;dino_sprite[2][51][69] = 1;dino_sprite[2][51][70] = 1;dino_sprite[2][51][71] = 1;dino_sprite[2][51][72] = 1;dino_sprite[2][51][73] = 1;dino_sprite[2][51][74] = 1;dino_sprite[2][51][75] = 1;dino_sprite[2][51][76] = 1;dino_sprite[2][51][77] = 1;dino_sprite[2][51][78] = 1;dino_sprite[2][51][79] = 1;dino_sprite[2][51][80] = 1;dino_sprite[2][51][81] = 1;dino_sprite[2][51][82] = 1;dino_sprite[2][51][83] = 1;dino_sprite[2][51][84] = 1;dino_sprite[2][51][85] = 1;dino_sprite[2][51][86] = 1;dino_sprite[2][51][87] = 1;dino_sprite[2][51][88] = 1;dino_sprite[2][51][89] = 1;dino_sprite[2][51][90] = 1;dino_sprite[2][51][91] = 1;dino_sprite[2][51][92] = 1;dino_sprite[2][52][3] = 1;dino_sprite[2][52][4] = 1;dino_sprite[2][52][5] = 1;dino_sprite[2][52][6] = 1;dino_sprite[2][52][7] = 1;dino_sprite[2][52][8] = 1;dino_sprite[2][52][9] = 1;dino_sprite[2][52][10] = 1;dino_sprite[2][52][11] = 1;dino_sprite[2][52][12] = 1;dino_sprite[2][52][13] = 1;dino_sprite[2][52][14] = 1;dino_sprite[2][52][15] = 1;dino_sprite[2][52][16] = 1;dino_sprite[2][52][17] = 1;dino_sprite[2][52][18] = 1;dino_sprite[2][52][19] = 1;dino_sprite[2][52][20] = 1;dino_sprite[2][52][21] = 1;dino_sprite[2][52][22] = 1;dino_sprite[2][52][23] = 1;dino_sprite[2][52][24] = 1;dino_sprite[2][52][25] = 1;dino_sprite[2][52][26] = 1;dino_sprite[2][52][27] = 1;dino_sprite[2][52][28] = 1;dino_sprite[2][52][29] = 1;dino_sprite[2][52][30] = 1;dino_sprite[2][52][31] = 1;dino_sprite[2][52][32] = 1;dino_sprite[2][52][33] = 1;dino_sprite[2][52][34] = 1;dino_sprite[2][52][35] = 1;dino_sprite[2][52][36] = 1;dino_sprite[2][52][37] = 1;dino_sprite[2][52][38] = 1;dino_sprite[2][52][39] = 1;dino_sprite[2][52][40] = 1;dino_sprite[2][52][41] = 1;dino_sprite[2][52][42] = 1;dino_sprite[2][52][43] = 1;dino_sprite[2][52][44] = 1;dino_sprite[2][52][45] = 1;dino_sprite[2][52][46] = 1;dino_sprite[2][52][47] = 1;dino_sprite[2][52][48] = 1;dino_sprite[2][52][49] = 1;dino_sprite[2][52][50] = 1;dino_sprite[2][52][51] = 1;dino_sprite[2][52][52] = 1;dino_sprite[2][52][53] = 1;dino_sprite[2][52][54] = 1;dino_sprite[2][52][55] = 1;dino_sprite[2][52][56] = 1;dino_sprite[2][52][57] = 1;dino_sprite[2][52][58] = 1;dino_sprite[2][52][59] = 1;dino_sprite[2][52][60] = 1;dino_sprite[2][52][61] = 1;dino_sprite[2][52][62] = 1;dino_sprite[2][52][63] = 1;dino_sprite[2][52][64] = 1;dino_sprite[2][52][65] = 1;dino_sprite[2][52][66] = 1;dino_sprite[2][52][67] = 1;dino_sprite[2][52][68] = 1;dino_sprite[2][52][69] = 1;dino_sprite[2][52][70] = 1;dino_sprite[2][52][71] = 1;dino_sprite[2][52][72] = 1;dino_sprite[2][52][73] = 1;dino_sprite[2][52][74] = 1;dino_sprite[2][52][75] = 1;dino_sprite[2][52][76] = 1;dino_sprite[2][52][77] = 1;dino_sprite[2][52][78] = 1;dino_sprite[2][52][79] = 1;dino_sprite[2][52][80] = 1;dino_sprite[2][52][81] = 1;dino_sprite[2][52][82] = 1;dino_sprite[2][52][83] = 1;dino_sprite[2][52][84] = 1;dino_sprite[2][52][85] = 1;dino_sprite[2][52][86] = 1;dino_sprite[2][52][87] = 1;dino_sprite[2][52][88] = 1;dino_sprite[2][52][89] = 1;dino_sprite[2][52][90] = 1;dino_sprite[2][52][91] = 1;dino_sprite[2][52][92] = 1;dino_sprite[2][53][3] = 1;dino_sprite[2][53][4] = 1;dino_sprite[2][53][5] = 1;dino_sprite[2][53][6] = 1;dino_sprite[2][53][7] = 1;dino_sprite[2][53][8] = 1;dino_sprite[2][53][9] = 1;dino_sprite[2][53][10] = 1;dino_sprite[2][53][11] = 1;dino_sprite[2][53][12] = 1;dino_sprite[2][53][13] = 1;dino_sprite[2][53][14] = 1;dino_sprite[2][53][15] = 1;dino_sprite[2][53][16] = 1;dino_sprite[2][53][17] = 1;dino_sprite[2][53][18] = 1;dino_sprite[2][53][19] = 1;dino_sprite[2][53][20] = 1;dino_sprite[2][53][21] = 1;dino_sprite[2][53][22] = 1;dino_sprite[2][53][23] = 1;dino_sprite[2][53][24] = 1;dino_sprite[2][53][25] = 1;dino_sprite[2][53][26] = 1;dino_sprite[2][53][27] = 1;dino_sprite[2][53][28] = 1;dino_sprite[2][53][29] = 1;dino_sprite[2][53][30] = 1;dino_sprite[2][53][31] = 1;dino_sprite[2][53][32] = 1;dino_sprite[2][53][33] = 1;dino_sprite[2][53][34] = 1;dino_sprite[2][53][35] = 1;dino_sprite[2][53][36] = 1;dino_sprite[2][53][37] = 1;dino_sprite[2][53][38] = 1;dino_sprite[2][53][39] = 1;dino_sprite[2][53][40] = 1;dino_sprite[2][53][41] = 1;dino_sprite[2][53][42] = 1;dino_sprite[2][53][43] = 1;dino_sprite[2][53][44] = 1;dino_sprite[2][53][45] = 1;dino_sprite[2][53][46] = 1;dino_sprite[2][53][47] = 1;dino_sprite[2][53][48] = 1;dino_sprite[2][53][49] = 1;dino_sprite[2][53][50] = 1;dino_sprite[2][53][51] = 1;dino_sprite[2][53][52] = 1;dino_sprite[2][53][53] = 1;dino_sprite[2][53][54] = 1;dino_sprite[2][53][55] = 1;dino_sprite[2][53][56] = 1;dino_sprite[2][53][57] = 1;dino_sprite[2][53][58] = 1;dino_sprite[2][53][59] = 1;dino_sprite[2][53][60] = 1;dino_sprite[2][53][61] = 1;dino_sprite[2][53][62] = 1;dino_sprite[2][53][63] = 1;dino_sprite[2][53][64] = 1;dino_sprite[2][53][65] = 1;dino_sprite[2][53][66] = 1;dino_sprite[2][53][67] = 1;dino_sprite[2][53][68] = 1;dino_sprite[2][53][69] = 1;dino_sprite[2][53][70] = 1;dino_sprite[2][53][71] = 1;dino_sprite[2][53][72] = 1;dino_sprite[2][53][73] = 1;dino_sprite[2][53][74] = 1;dino_sprite[2][53][75] = 1;dino_sprite[2][53][76] = 1;dino_sprite[2][53][77] = 1;dino_sprite[2][53][78] = 1;dino_sprite[2][53][79] = 1;dino_sprite[2][53][80] = 1;dino_sprite[2][53][81] = 1;dino_sprite[2][53][82] = 1;dino_sprite[2][53][83] = 1;dino_sprite[2][53][84] = 1;dino_sprite[2][53][85] = 1;dino_sprite[2][53][86] = 1;dino_sprite[2][53][87] = 1;dino_sprite[2][53][88] = 1;dino_sprite[2][53][89] = 1;dino_sprite[2][53][90] = 1;dino_sprite[2][53][91] = 1;dino_sprite[2][53][92] = 1;dino_sprite[2][54][3] = 1;dino_sprite[2][54][4] = 1;dino_sprite[2][54][5] = 1;dino_sprite[2][54][6] = 1;dino_sprite[2][54][7] = 1;dino_sprite[2][54][8] = 1;dino_sprite[2][54][9] = 1;dino_sprite[2][54][10] = 1;dino_sprite[2][54][11] = 1;dino_sprite[2][54][12] = 1;dino_sprite[2][54][13] = 1;dino_sprite[2][54][14] = 1;dino_sprite[2][54][15] = 1;dino_sprite[2][54][16] = 1;dino_sprite[2][54][17] = 1;dino_sprite[2][54][18] = 1;dino_sprite[2][54][19] = 1;dino_sprite[2][54][20] = 1;dino_sprite[2][54][21] = 1;dino_sprite[2][54][22] = 1;dino_sprite[2][54][23] = 1;dino_sprite[2][54][24] = 1;dino_sprite[2][54][25] = 1;dino_sprite[2][54][26] = 1;dino_sprite[2][54][27] = 1;dino_sprite[2][54][28] = 1;dino_sprite[2][54][29] = 1;dino_sprite[2][54][30] = 1;dino_sprite[2][54][31] = 1;dino_sprite[2][54][32] = 1;dino_sprite[2][54][33] = 1;dino_sprite[2][54][34] = 1;dino_sprite[2][54][35] = 1;dino_sprite[2][54][36] = 1;dino_sprite[2][54][37] = 1;dino_sprite[2][54][38] = 1;dino_sprite[2][54][39] = 1;dino_sprite[2][54][40] = 1;dino_sprite[2][54][41] = 1;dino_sprite[2][54][42] = 1;dino_sprite[2][54][43] = 1;dino_sprite[2][54][44] = 1;dino_sprite[2][54][45] = 1;dino_sprite[2][54][46] = 1;dino_sprite[2][54][47] = 1;dino_sprite[2][54][48] = 1;dino_sprite[2][54][49] = 1;dino_sprite[2][54][50] = 1;dino_sprite[2][54][51] = 1;dino_sprite[2][54][52] = 1;dino_sprite[2][54][53] = 1;dino_sprite[2][54][54] = 1;dino_sprite[2][54][55] = 1;dino_sprite[2][54][56] = 1;dino_sprite[2][54][57] = 1;dino_sprite[2][54][58] = 1;dino_sprite[2][54][59] = 1;dino_sprite[2][54][60] = 1;dino_sprite[2][54][61] = 1;dino_sprite[2][54][62] = 1;dino_sprite[2][54][63] = 1;dino_sprite[2][54][64] = 1;dino_sprite[2][54][65] = 1;dino_sprite[2][54][66] = 1;dino_sprite[2][54][67] = 1;dino_sprite[2][54][68] = 1;dino_sprite[2][54][69] = 1;dino_sprite[2][54][70] = 1;dino_sprite[2][54][71] = 1;dino_sprite[2][54][72] = 1;dino_sprite[2][54][73] = 1;dino_sprite[2][54][74] = 1;dino_sprite[2][54][75] = 1;dino_sprite[2][54][76] = 1;dino_sprite[2][54][77] = 1;dino_sprite[2][54][78] = 1;dino_sprite[2][54][79] = 1;dino_sprite[2][54][80] = 1;dino_sprite[2][54][81] = 1;dino_sprite[2][54][82] = 1;dino_sprite[2][54][83] = 1;dino_sprite[2][54][84] = 1;dino_sprite[2][54][85] = 1;dino_sprite[2][54][86] = 1;dino_sprite[2][54][87] = 1;dino_sprite[2][54][88] = 1;dino_sprite[2][54][89] = 1;dino_sprite[2][54][90] = 1;dino_sprite[2][54][91] = 1;dino_sprite[2][54][92] = 1;dino_sprite[2][55][3] = 1;dino_sprite[2][55][4] = 1;dino_sprite[2][55][5] = 1;dino_sprite[2][55][6] = 1;dino_sprite[2][55][7] = 1;dino_sprite[2][55][8] = 1;dino_sprite[2][55][9] = 1;dino_sprite[2][55][10] = 1;dino_sprite[2][55][11] = 1;dino_sprite[2][55][12] = 1;dino_sprite[2][55][13] = 1;dino_sprite[2][55][14] = 1;dino_sprite[2][55][15] = 1;dino_sprite[2][55][16] = 1;dino_sprite[2][55][17] = 1;dino_sprite[2][55][18] = 1;dino_sprite[2][55][19] = 1;dino_sprite[2][55][20] = 1;dino_sprite[2][55][21] = 1;dino_sprite[2][55][22] = 1;dino_sprite[2][55][23] = 1;dino_sprite[2][55][24] = 1;dino_sprite[2][55][25] = 1;dino_sprite[2][55][26] = 1;dino_sprite[2][55][27] = 1;dino_sprite[2][55][28] = 1;dino_sprite[2][55][29] = 1;dino_sprite[2][55][30] = 1;dino_sprite[2][55][31] = 1;dino_sprite[2][55][32] = 1;dino_sprite[2][55][33] = 1;dino_sprite[2][55][34] = 1;dino_sprite[2][55][35] = 1;dino_sprite[2][55][36] = 1;dino_sprite[2][55][37] = 1;dino_sprite[2][55][38] = 1;dino_sprite[2][55][39] = 1;dino_sprite[2][55][40] = 1;dino_sprite[2][55][41] = 1;dino_sprite[2][55][42] = 1;dino_sprite[2][55][43] = 1;dino_sprite[2][55][44] = 1;dino_sprite[2][55][45] = 1;dino_sprite[2][55][46] = 1;dino_sprite[2][55][47] = 1;dino_sprite[2][55][48] = 1;dino_sprite[2][55][49] = 1;dino_sprite[2][55][50] = 1;dino_sprite[2][55][51] = 1;dino_sprite[2][55][52] = 1;dino_sprite[2][55][53] = 1;dino_sprite[2][55][54] = 1;dino_sprite[2][55][55] = 1;dino_sprite[2][55][56] = 1;dino_sprite[2][55][57] = 1;dino_sprite[2][55][58] = 1;dino_sprite[2][55][59] = 1;dino_sprite[2][55][60] = 1;dino_sprite[2][55][61] = 1;dino_sprite[2][55][62] = 1;dino_sprite[2][55][63] = 1;dino_sprite[2][55][64] = 1;dino_sprite[2][55][65] = 1;dino_sprite[2][55][66] = 1;dino_sprite[2][55][67] = 1;dino_sprite[2][55][68] = 1;dino_sprite[2][55][69] = 1;dino_sprite[2][55][70] = 1;dino_sprite[2][55][71] = 1;dino_sprite[2][55][72] = 1;dino_sprite[2][55][73] = 1;dino_sprite[2][55][74] = 1;dino_sprite[2][55][75] = 1;dino_sprite[2][55][76] = 1;dino_sprite[2][55][77] = 1;dino_sprite[2][55][78] = 1;dino_sprite[2][55][79] = 1;dino_sprite[2][55][80] = 1;dino_sprite[2][55][81] = 1;dino_sprite[2][55][82] = 1;dino_sprite[2][55][83] = 1;dino_sprite[2][55][84] = 1;dino_sprite[2][55][85] = 1;dino_sprite[2][55][86] = 1;dino_sprite[2][55][87] = 1;dino_sprite[2][55][88] = 1;dino_sprite[2][55][89] = 1;dino_sprite[2][55][90] = 1;dino_sprite[2][55][91] = 1;dino_sprite[2][55][92] = 1;dino_sprite[2][56][0] = 1;dino_sprite[2][56][1] = 1;dino_sprite[2][56][2] = 1;dino_sprite[2][56][3] = 1;dino_sprite[2][56][4] = 1;dino_sprite[2][56][5] = 1;dino_sprite[2][56][6] = 1;dino_sprite[2][56][7] = 1;dino_sprite[2][56][8] = 1;dino_sprite[2][56][9] = 1;dino_sprite[2][56][10] = 1;dino_sprite[2][56][11] = 1;dino_sprite[2][56][12] = 1;dino_sprite[2][56][13] = 1;dino_sprite[2][56][14] = 1;dino_sprite[2][56][15] = 1;dino_sprite[2][56][16] = 1;dino_sprite[2][56][17] = 1;dino_sprite[2][56][18] = 1;dino_sprite[2][56][19] = 1;dino_sprite[2][56][20] = 1;dino_sprite[2][56][21] = 1;dino_sprite[2][56][22] = 1;dino_sprite[2][56][23] = 1;dino_sprite[2][56][24] = 1;dino_sprite[2][56][25] = 1;dino_sprite[2][56][26] = 1;dino_sprite[2][56][27] = 1;dino_sprite[2][56][28] = 1;dino_sprite[2][56][29] = 1;dino_sprite[2][56][30] = 1;dino_sprite[2][56][31] = 1;dino_sprite[2][56][32] = 1;dino_sprite[2][56][33] = 1;dino_sprite[2][56][34] = 1;dino_sprite[2][56][35] = 1;dino_sprite[2][56][36] = 1;dino_sprite[2][56][37] = 1;dino_sprite[2][56][38] = 1;dino_sprite[2][56][39] = 1;dino_sprite[2][56][40] = 1;dino_sprite[2][56][41] = 1;dino_sprite[2][56][42] = 1;dino_sprite[2][56][43] = 1;dino_sprite[2][56][44] = 1;dino_sprite[2][56][45] = 1;dino_sprite[2][56][46] = 1;dino_sprite[2][56][47] = 1;dino_sprite[2][56][48] = 1;dino_sprite[2][56][49] = 1;dino_sprite[2][56][50] = 1;dino_sprite[2][56][51] = 1;dino_sprite[2][56][52] = 1;dino_sprite[2][56][53] = 1;dino_sprite[2][56][54] = 1;dino_sprite[2][56][55] = 1;dino_sprite[2][56][56] = 1;dino_sprite[2][56][57] = 1;dino_sprite[2][56][58] = 1;dino_sprite[2][56][59] = 1;dino_sprite[2][56][60] = 1;dino_sprite[2][56][61] = 1;dino_sprite[2][56][62] = 1;dino_sprite[2][56][63] = 1;dino_sprite[2][56][64] = 1;dino_sprite[2][56][65] = 1;dino_sprite[2][56][66] = 1;dino_sprite[2][56][67] = 1;dino_sprite[2][56][68] = 1;dino_sprite[2][56][69] = 1;dino_sprite[2][56][70] = 1;dino_sprite[2][56][71] = 1;dino_sprite[2][56][72] = 1;dino_sprite[2][56][73] = 1;dino_sprite[2][56][74] = 1;dino_sprite[2][56][75] = 1;dino_sprite[2][56][76] = 1;dino_sprite[2][56][77] = 1;dino_sprite[2][56][89] = 1;dino_sprite[2][56][90] = 1;dino_sprite[2][56][91] = 1;dino_sprite[2][56][92] = 1;dino_sprite[2][57][0] = 1;dino_sprite[2][57][1] = 1;dino_sprite[2][57][2] = 1;dino_sprite[2][57][3] = 1;dino_sprite[2][57][4] = 1;dino_sprite[2][57][5] = 1;dino_sprite[2][57][6] = 1;dino_sprite[2][57][7] = 1;dino_sprite[2][57][8] = 1;dino_sprite[2][57][9] = 1;dino_sprite[2][57][10] = 1;dino_sprite[2][57][11] = 1;dino_sprite[2][57][12] = 1;dino_sprite[2][57][13] = 1;dino_sprite[2][57][14] = 1;dino_sprite[2][57][15] = 1;dino_sprite[2][57][16] = 1;dino_sprite[2][57][17] = 1;dino_sprite[2][57][18] = 1;dino_sprite[2][57][19] = 1;dino_sprite[2][57][20] = 1;dino_sprite[2][57][21] = 1;dino_sprite[2][57][22] = 1;dino_sprite[2][57][23] = 1;dino_sprite[2][57][24] = 1;dino_sprite[2][57][25] = 1;dino_sprite[2][57][26] = 1;dino_sprite[2][57][27] = 1;dino_sprite[2][57][28] = 1;dino_sprite[2][57][29] = 1;dino_sprite[2][57][30] = 1;dino_sprite[2][57][31] = 1;dino_sprite[2][57][32] = 1;dino_sprite[2][57][33] = 1;dino_sprite[2][57][34] = 1;dino_sprite[2][57][35] = 1;dino_sprite[2][57][36] = 1;dino_sprite[2][57][37] = 1;dino_sprite[2][57][38] = 1;dino_sprite[2][57][39] = 1;dino_sprite[2][57][40] = 1;dino_sprite[2][57][41] = 1;dino_sprite[2][57][42] = 1;dino_sprite[2][57][43] = 1;dino_sprite[2][57][44] = 1;dino_sprite[2][57][45] = 1;dino_sprite[2][57][46] = 1;dino_sprite[2][57][47] = 1;dino_sprite[2][57][48] = 1;dino_sprite[2][57][49] = 1;dino_sprite[2][57][50] = 1;dino_sprite[2][57][51] = 1;dino_sprite[2][57][52] = 1;dino_sprite[2][57][53] = 1;dino_sprite[2][57][54] = 1;dino_sprite[2][57][55] = 1;dino_sprite[2][57][56] = 1;dino_sprite[2][57][57] = 1;dino_sprite[2][57][58] = 1;dino_sprite[2][57][59] = 1;dino_sprite[2][57][60] = 1;dino_sprite[2][57][61] = 1;dino_sprite[2][57][62] = 1;dino_sprite[2][57][63] = 1;dino_sprite[2][57][64] = 1;dino_sprite[2][57][65] = 1;dino_sprite[2][57][66] = 1;dino_sprite[2][57][67] = 1;dino_sprite[2][57][68] = 1;dino_sprite[2][57][69] = 1;dino_sprite[2][57][70] = 1;dino_sprite[2][57][71] = 1;dino_sprite[2][57][72] = 1;dino_sprite[2][57][73] = 1;dino_sprite[2][57][74] = 1;dino_sprite[2][57][75] = 1;dino_sprite[2][57][76] = 1;dino_sprite[2][57][77] = 1;dino_sprite[2][57][89] = 1;dino_sprite[2][57][90] = 1;dino_sprite[2][57][91] = 1;dino_sprite[2][57][92] = 1;dino_sprite[2][58][0] = 1;dino_sprite[2][58][1] = 1;dino_sprite[2][58][2] = 1;dino_sprite[2][58][3] = 1;dino_sprite[2][58][4] = 1;dino_sprite[2][58][5] = 1;dino_sprite[2][58][6] = 1;dino_sprite[2][58][7] = 1;dino_sprite[2][58][8] = 1;dino_sprite[2][58][9] = 1;dino_sprite[2][58][10] = 1;dino_sprite[2][58][11] = 1;dino_sprite[2][58][12] = 1;dino_sprite[2][58][13] = 1;dino_sprite[2][58][14] = 1;dino_sprite[2][58][15] = 1;dino_sprite[2][58][16] = 1;dino_sprite[2][58][17] = 1;dino_sprite[2][58][18] = 1;dino_sprite[2][58][19] = 1;dino_sprite[2][58][20] = 1;dino_sprite[2][58][21] = 1;dino_sprite[2][58][22] = 1;dino_sprite[2][58][23] = 1;dino_sprite[2][58][24] = 1;dino_sprite[2][58][25] = 1;dino_sprite[2][58][26] = 1;dino_sprite[2][58][27] = 1;dino_sprite[2][58][28] = 1;dino_sprite[2][58][29] = 1;dino_sprite[2][58][30] = 1;dino_sprite[2][58][31] = 1;dino_sprite[2][58][32] = 1;dino_sprite[2][58][33] = 1;dino_sprite[2][58][34] = 1;dino_sprite[2][58][35] = 1;dino_sprite[2][58][36] = 1;dino_sprite[2][58][37] = 1;dino_sprite[2][58][38] = 1;dino_sprite[2][58][39] = 1;dino_sprite[2][58][40] = 1;dino_sprite[2][58][41] = 1;dino_sprite[2][58][42] = 1;dino_sprite[2][58][43] = 1;dino_sprite[2][58][44] = 1;dino_sprite[2][58][45] = 1;dino_sprite[2][58][46] = 1;dino_sprite[2][58][47] = 1;dino_sprite[2][58][48] = 1;dino_sprite[2][58][49] = 1;dino_sprite[2][58][50] = 1;dino_sprite[2][58][51] = 1;dino_sprite[2][58][52] = 1;dino_sprite[2][58][53] = 1;dino_sprite[2][58][54] = 1;dino_sprite[2][58][55] = 1;dino_sprite[2][58][56] = 1;dino_sprite[2][58][57] = 1;dino_sprite[2][58][58] = 1;dino_sprite[2][58][59] = 1;dino_sprite[2][58][60] = 1;dino_sprite[2][58][61] = 1;dino_sprite[2][58][62] = 1;dino_sprite[2][58][63] = 1;dino_sprite[2][58][64] = 1;dino_sprite[2][58][65] = 1;dino_sprite[2][58][66] = 1;dino_sprite[2][58][67] = 1;dino_sprite[2][58][68] = 1;dino_sprite[2][58][69] = 1;dino_sprite[2][58][70] = 1;dino_sprite[2][58][71] = 1;dino_sprite[2][58][72] = 1;dino_sprite[2][58][73] = 1;dino_sprite[2][58][74] = 1;dino_sprite[2][58][75] = 1;dino_sprite[2][58][76] = 1;dino_sprite[2][58][77] = 1;dino_sprite[2][58][89] = 1;dino_sprite[2][58][90] = 1;dino_sprite[2][58][91] = 1;dino_sprite[2][58][92] = 1;dino_sprite[2][58][95] = 1;dino_sprite[2][59][0] = 1;dino_sprite[2][59][1] = 1;dino_sprite[2][59][2] = 1;dino_sprite[2][59][3] = 1;dino_sprite[2][59][4] = 1;dino_sprite[2][59][5] = 1;dino_sprite[2][59][6] = 1;dino_sprite[2][59][7] = 1;dino_sprite[2][59][8] = 1;dino_sprite[2][59][9] = 1;dino_sprite[2][59][10] = 1;dino_sprite[2][59][11] = 1;dino_sprite[2][59][12] = 1;dino_sprite[2][59][13] = 1;dino_sprite[2][59][14] = 1;dino_sprite[2][59][15] = 1;dino_sprite[2][59][16] = 1;dino_sprite[2][59][17] = 1;dino_sprite[2][59][18] = 1;dino_sprite[2][59][19] = 1;dino_sprite[2][59][20] = 1;dino_sprite[2][59][21] = 1;dino_sprite[2][59][22] = 1;dino_sprite[2][59][23] = 1;dino_sprite[2][59][24] = 1;dino_sprite[2][59][25] = 1;dino_sprite[2][59][26] = 1;dino_sprite[2][59][27] = 1;dino_sprite[2][59][28] = 1;dino_sprite[2][59][29] = 1;dino_sprite[2][59][30] = 1;dino_sprite[2][59][31] = 1;dino_sprite[2][59][32] = 1;dino_sprite[2][59][33] = 1;dino_sprite[2][59][34] = 1;dino_sprite[2][59][35] = 1;dino_sprite[2][59][36] = 1;dino_sprite[2][59][37] = 1;dino_sprite[2][59][38] = 1;dino_sprite[2][59][39] = 1;dino_sprite[2][59][40] = 1;dino_sprite[2][59][41] = 1;dino_sprite[2][59][42] = 1;dino_sprite[2][59][43] = 1;dino_sprite[2][59][44] = 1;dino_sprite[2][59][45] = 1;dino_sprite[2][59][46] = 1;dino_sprite[2][59][47] = 1;dino_sprite[2][59][48] = 1;dino_sprite[2][59][49] = 1;dino_sprite[2][59][50] = 1;dino_sprite[2][59][51] = 1;dino_sprite[2][59][52] = 1;dino_sprite[2][59][53] = 1;dino_sprite[2][59][54] = 1;dino_sprite[2][59][55] = 1;dino_sprite[2][59][56] = 1;dino_sprite[2][59][57] = 1;dino_sprite[2][59][58] = 1;dino_sprite[2][59][59] = 1;dino_sprite[2][59][60] = 1;dino_sprite[2][59][61] = 1;dino_sprite[2][59][62] = 1;dino_sprite[2][59][63] = 1;dino_sprite[2][59][64] = 1;dino_sprite[2][59][65] = 1;dino_sprite[2][59][66] = 1;dino_sprite[2][59][67] = 1;dino_sprite[2][59][68] = 1;dino_sprite[2][59][69] = 1;dino_sprite[2][59][70] = 1;dino_sprite[2][59][71] = 1;dino_sprite[2][59][72] = 1;dino_sprite[2][59][73] = 1;dino_sprite[2][59][74] = 1;dino_sprite[2][59][75] = 1;dino_sprite[2][59][76] = 1;dino_sprite[2][59][77] = 1;dino_sprite[2][59][89] = 1;dino_sprite[2][59][90] = 1;dino_sprite[2][59][91] = 1;dino_sprite[2][59][92] = 1;dino_sprite[2][59][95] = 1;dino_sprite[2][60][0] = 1;dino_sprite[2][60][1] = 1;dino_sprite[2][60][2] = 1;dino_sprite[2][60][3] = 1;dino_sprite[2][60][4] = 1;dino_sprite[2][60][5] = 1;dino_sprite[2][60][6] = 1;dino_sprite[2][60][7] = 1;dino_sprite[2][60][8] = 1;dino_sprite[2][60][9] = 1;dino_sprite[2][60][10] = 1;dino_sprite[2][60][11] = 1;dino_sprite[2][60][12] = 1;dino_sprite[2][60][13] = 1;dino_sprite[2][60][14] = 1;dino_sprite[2][60][15] = 1;dino_sprite[2][60][16] = 1;dino_sprite[2][60][17] = 1;dino_sprite[2][60][18] = 1;dino_sprite[2][60][19] = 1;dino_sprite[2][60][20] = 1;dino_sprite[2][60][21] = 1;dino_sprite[2][60][22] = 1;dino_sprite[2][60][23] = 1;dino_sprite[2][60][24] = 1;dino_sprite[2][60][25] = 1;dino_sprite[2][60][26] = 1;dino_sprite[2][60][27] = 1;dino_sprite[2][60][28] = 1;dino_sprite[2][60][29] = 1;dino_sprite[2][60][30] = 1;dino_sprite[2][60][31] = 1;dino_sprite[2][60][32] = 1;dino_sprite[2][60][33] = 1;dino_sprite[2][60][34] = 1;dino_sprite[2][60][35] = 1;dino_sprite[2][60][36] = 1;dino_sprite[2][60][37] = 1;dino_sprite[2][60][38] = 1;dino_sprite[2][60][39] = 1;dino_sprite[2][60][40] = 1;dino_sprite[2][60][41] = 1;dino_sprite[2][60][42] = 1;dino_sprite[2][60][43] = 1;dino_sprite[2][60][44] = 1;dino_sprite[2][60][45] = 1;dino_sprite[2][60][46] = 1;dino_sprite[2][60][47] = 1;dino_sprite[2][60][48] = 1;dino_sprite[2][60][49] = 1;dino_sprite[2][60][50] = 1;dino_sprite[2][60][51] = 1;dino_sprite[2][60][52] = 1;dino_sprite[2][60][53] = 1;dino_sprite[2][60][54] = 1;dino_sprite[2][60][55] = 1;dino_sprite[2][60][56] = 1;dino_sprite[2][60][57] = 1;dino_sprite[2][60][58] = 1;dino_sprite[2][60][59] = 1;dino_sprite[2][60][60] = 1;dino_sprite[2][60][61] = 1;dino_sprite[2][60][62] = 1;dino_sprite[2][60][63] = 1;dino_sprite[2][60][64] = 1;dino_sprite[2][60][65] = 1;dino_sprite[2][60][66] = 1;dino_sprite[2][60][67] = 1;dino_sprite[2][60][68] = 1;dino_sprite[2][60][69] = 1;dino_sprite[2][60][70] = 1;dino_sprite[2][60][71] = 1;dino_sprite[2][60][72] = 1;dino_sprite[2][60][73] = 1;dino_sprite[2][60][74] = 1;dino_sprite[2][60][75] = 1;dino_sprite[2][60][76] = 1;dino_sprite[2][60][77] = 1;dino_sprite[2][60][89] = 1;dino_sprite[2][60][90] = 1;dino_sprite[2][60][91] = 1;dino_sprite[2][60][92] = 1;dino_sprite[2][61][0] = 1;dino_sprite[2][61][1] = 1;dino_sprite[2][61][2] = 1;dino_sprite[2][61][3] = 1;dino_sprite[2][61][4] = 1;dino_sprite[2][61][5] = 1;dino_sprite[2][61][6] = 1;dino_sprite[2][61][10] = 1;dino_sprite[2][61][11] = 1;dino_sprite[2][61][12] = 1;dino_sprite[2][61][13] = 1;dino_sprite[2][61][14] = 1;dino_sprite[2][61][15] = 1;dino_sprite[2][61][16] = 1;dino_sprite[2][61][17] = 1;dino_sprite[2][61][18] = 1;dino_sprite[2][61][19] = 1;dino_sprite[2][61][20] = 1;dino_sprite[2][61][21] = 1;dino_sprite[2][61][22] = 1;dino_sprite[2][61][23] = 1;dino_sprite[2][61][24] = 1;dino_sprite[2][61][25] = 1;dino_sprite[2][61][26] = 1;dino_sprite[2][61][27] = 1;dino_sprite[2][61][28] = 1;dino_sprite[2][61][29] = 1;dino_sprite[2][61][30] = 1;dino_sprite[2][61][31] = 1;dino_sprite[2][61][32] = 1;dino_sprite[2][61][33] = 1;dino_sprite[2][61][34] = 1;dino_sprite[2][61][35] = 1;dino_sprite[2][61][36] = 1;dino_sprite[2][61][37] = 1;dino_sprite[2][61][38] = 1;dino_sprite[2][61][39] = 1;dino_sprite[2][61][40] = 1;dino_sprite[2][61][41] = 1;dino_sprite[2][61][42] = 1;dino_sprite[2][61][43] = 1;dino_sprite[2][61][44] = 1;dino_sprite[2][61][45] = 1;dino_sprite[2][61][46] = 1;dino_sprite[2][61][47] = 1;dino_sprite[2][61][48] = 1;dino_sprite[2][61][49] = 1;dino_sprite[2][61][50] = 1;dino_sprite[2][61][51] = 1;dino_sprite[2][61][52] = 1;dino_sprite[2][61][53] = 1;dino_sprite[2][61][54] = 1;dino_sprite[2][61][55] = 1;dino_sprite[2][61][56] = 1;dino_sprite[2][61][57] = 1;dino_sprite[2][61][58] = 1;dino_sprite[2][61][59] = 1;dino_sprite[2][61][60] = 1;dino_sprite[2][61][61] = 1;dino_sprite[2][61][62] = 1;dino_sprite[2][61][63] = 1;dino_sprite[2][61][64] = 1;dino_sprite[2][61][65] = 1;dino_sprite[2][61][66] = 1;dino_sprite[2][61][67] = 1;dino_sprite[2][61][68] = 1;dino_sprite[2][61][69] = 1;dino_sprite[2][61][70] = 1;dino_sprite[2][61][71] = 1;dino_sprite[2][61][72] = 1;dino_sprite[2][62][0] = 1;dino_sprite[2][62][1] = 1;dino_sprite[2][62][2] = 1;dino_sprite[2][62][3] = 1;dino_sprite[2][62][4] = 1;dino_sprite[2][62][5] = 1;dino_sprite[2][62][6] = 1;dino_sprite[2][62][10] = 1;dino_sprite[2][62][11] = 1;dino_sprite[2][62][12] = 1;dino_sprite[2][62][13] = 1;dino_sprite[2][62][14] = 1;dino_sprite[2][62][15] = 1;dino_sprite[2][62][16] = 1;dino_sprite[2][62][17] = 1;dino_sprite[2][62][18] = 1;dino_sprite[2][62][19] = 1;dino_sprite[2][62][20] = 1;dino_sprite[2][62][21] = 1;dino_sprite[2][62][22] = 1;dino_sprite[2][62][23] = 1;dino_sprite[2][62][24] = 1;dino_sprite[2][62][25] = 1;dino_sprite[2][62][26] = 1;dino_sprite[2][62][27] = 1;dino_sprite[2][62][28] = 1;dino_sprite[2][62][29] = 1;dino_sprite[2][62][30] = 1;dino_sprite[2][62][31] = 1;dino_sprite[2][62][32] = 1;dino_sprite[2][62][33] = 1;dino_sprite[2][62][34] = 1;dino_sprite[2][62][35] = 1;dino_sprite[2][62][36] = 1;dino_sprite[2][62][37] = 1;dino_sprite[2][62][38] = 1;dino_sprite[2][62][39] = 1;dino_sprite[2][62][40] = 1;dino_sprite[2][62][41] = 1;dino_sprite[2][62][42] = 1;dino_sprite[2][62][43] = 1;dino_sprite[2][62][44] = 1;dino_sprite[2][62][45] = 1;dino_sprite[2][62][46] = 1;dino_sprite[2][62][47] = 1;dino_sprite[2][62][48] = 1;dino_sprite[2][62][49] = 1;dino_sprite[2][62][50] = 1;dino_sprite[2][62][51] = 1;dino_sprite[2][62][52] = 1;dino_sprite[2][62][53] = 1;dino_sprite[2][62][54] = 1;dino_sprite[2][62][55] = 1;dino_sprite[2][62][56] = 1;dino_sprite[2][62][57] = 1;dino_sprite[2][62][58] = 1;dino_sprite[2][62][59] = 1;dino_sprite[2][62][60] = 1;dino_sprite[2][62][61] = 1;dino_sprite[2][62][62] = 1;dino_sprite[2][62][63] = 1;dino_sprite[2][62][64] = 1;dino_sprite[2][62][65] = 1;dino_sprite[2][62][66] = 1;dino_sprite[2][62][67] = 1;dino_sprite[2][62][68] = 1;dino_sprite[2][62][69] = 1;dino_sprite[2][62][70] = 1;dino_sprite[2][62][71] = 1;dino_sprite[2][62][72] = 1;dino_sprite[2][63][0] = 1;dino_sprite[2][63][1] = 1;dino_sprite[2][63][2] = 1;dino_sprite[2][63][3] = 1;dino_sprite[2][63][4] = 1;dino_sprite[2][63][5] = 1;dino_sprite[2][63][6] = 1;dino_sprite[2][63][10] = 1;dino_sprite[2][63][11] = 1;dino_sprite[2][63][12] = 1;dino_sprite[2][63][13] = 1;dino_sprite[2][63][14] = 1;dino_sprite[2][63][15] = 1;dino_sprite[2][63][16] = 1;dino_sprite[2][63][17] = 1;dino_sprite[2][63][18] = 1;dino_sprite[2][63][19] = 1;dino_sprite[2][63][20] = 1;dino_sprite[2][63][21] = 1;dino_sprite[2][63][22] = 1;dino_sprite[2][63][23] = 1;dino_sprite[2][63][24] = 1;dino_sprite[2][63][25] = 1;dino_sprite[2][63][26] = 1;dino_sprite[2][63][27] = 1;dino_sprite[2][63][28] = 1;dino_sprite[2][63][29] = 1;dino_sprite[2][63][30] = 1;dino_sprite[2][63][31] = 1;dino_sprite[2][63][32] = 1;dino_sprite[2][63][33] = 1;dino_sprite[2][63][34] = 1;dino_sprite[2][63][35] = 1;dino_sprite[2][63][36] = 1;dino_sprite[2][63][37] = 1;dino_sprite[2][63][38] = 1;dino_sprite[2][63][39] = 1;dino_sprite[2][63][40] = 1;dino_sprite[2][63][41] = 1;dino_sprite[2][63][42] = 1;dino_sprite[2][63][43] = 1;dino_sprite[2][63][44] = 1;dino_sprite[2][63][45] = 1;dino_sprite[2][63][46] = 1;dino_sprite[2][63][47] = 1;dino_sprite[2][63][48] = 1;dino_sprite[2][63][49] = 1;dino_sprite[2][63][50] = 1;dino_sprite[2][63][51] = 1;dino_sprite[2][63][52] = 1;dino_sprite[2][63][53] = 1;dino_sprite[2][63][54] = 1;dino_sprite[2][63][55] = 1;dino_sprite[2][63][56] = 1;dino_sprite[2][63][57] = 1;dino_sprite[2][63][58] = 1;dino_sprite[2][63][59] = 1;dino_sprite[2][63][60] = 1;dino_sprite[2][63][61] = 1;dino_sprite[2][63][62] = 1;dino_sprite[2][63][63] = 1;dino_sprite[2][63][64] = 1;dino_sprite[2][63][65] = 1;dino_sprite[2][63][66] = 1;dino_sprite[2][63][67] = 1;dino_sprite[2][63][68] = 1;dino_sprite[2][63][69] = 1;dino_sprite[2][63][70] = 1;dino_sprite[2][63][71] = 1;dino_sprite[2][63][72] = 1;dino_sprite[2][64][0] = 1;dino_sprite[2][64][1] = 1;dino_sprite[2][64][2] = 1;dino_sprite[2][64][3] = 1;dino_sprite[2][64][4] = 1;dino_sprite[2][64][5] = 1;dino_sprite[2][64][6] = 1;dino_sprite[2][64][10] = 1;dino_sprite[2][64][11] = 1;dino_sprite[2][64][12] = 1;dino_sprite[2][64][13] = 1;dino_sprite[2][64][14] = 1;dino_sprite[2][64][15] = 1;dino_sprite[2][64][16] = 1;dino_sprite[2][64][17] = 1;dino_sprite[2][64][18] = 1;dino_sprite[2][64][19] = 1;dino_sprite[2][64][20] = 1;dino_sprite[2][64][21] = 1;dino_sprite[2][64][22] = 1;dino_sprite[2][64][23] = 1;dino_sprite[2][64][24] = 1;dino_sprite[2][64][25] = 1;dino_sprite[2][64][26] = 1;dino_sprite[2][64][27] = 1;dino_sprite[2][64][28] = 1;dino_sprite[2][64][29] = 1;dino_sprite[2][64][30] = 1;dino_sprite[2][64][31] = 1;dino_sprite[2][64][32] = 1;dino_sprite[2][64][33] = 1;dino_sprite[2][64][34] = 1;dino_sprite[2][64][35] = 1;dino_sprite[2][64][36] = 1;dino_sprite[2][64][37] = 1;dino_sprite[2][64][38] = 1;dino_sprite[2][64][39] = 1;dino_sprite[2][64][40] = 1;dino_sprite[2][64][41] = 1;dino_sprite[2][64][42] = 1;dino_sprite[2][64][43] = 1;dino_sprite[2][64][44] = 1;dino_sprite[2][64][45] = 1;dino_sprite[2][64][46] = 1;dino_sprite[2][64][47] = 1;dino_sprite[2][64][48] = 1;dino_sprite[2][64][49] = 1;dino_sprite[2][64][50] = 1;dino_sprite[2][64][51] = 1;dino_sprite[2][64][52] = 1;dino_sprite[2][64][53] = 1;dino_sprite[2][64][54] = 1;dino_sprite[2][64][55] = 1;dino_sprite[2][64][56] = 1;dino_sprite[2][64][57] = 1;dino_sprite[2][64][58] = 1;dino_sprite[2][64][59] = 1;dino_sprite[2][64][60] = 1;dino_sprite[2][64][61] = 1;dino_sprite[2][64][62] = 1;dino_sprite[2][64][63] = 1;dino_sprite[2][64][64] = 1;dino_sprite[2][64][65] = 1;dino_sprite[2][64][66] = 1;dino_sprite[2][64][67] = 1;dino_sprite[2][64][68] = 1;dino_sprite[2][64][69] = 1;dino_sprite[2][64][70] = 1;dino_sprite[2][64][71] = 1;dino_sprite[2][64][72] = 1;dino_sprite[2][65][0] = 1;dino_sprite[2][65][1] = 1;dino_sprite[2][65][2] = 1;dino_sprite[2][65][3] = 1;dino_sprite[2][65][4] = 1;dino_sprite[2][65][5] = 1;dino_sprite[2][65][6] = 1;dino_sprite[2][65][8] = 1;dino_sprite[2][65][10] = 1;dino_sprite[2][65][11] = 1;dino_sprite[2][65][12] = 1;dino_sprite[2][65][13] = 1;dino_sprite[2][65][14] = 1;dino_sprite[2][65][15] = 1;dino_sprite[2][65][16] = 1;dino_sprite[2][65][17] = 1;dino_sprite[2][65][18] = 1;dino_sprite[2][65][19] = 1;dino_sprite[2][65][20] = 1;dino_sprite[2][65][21] = 1;dino_sprite[2][65][22] = 1;dino_sprite[2][65][23] = 1;dino_sprite[2][65][24] = 1;dino_sprite[2][65][25] = 1;dino_sprite[2][65][26] = 1;dino_sprite[2][65][27] = 1;dino_sprite[2][65][28] = 1;dino_sprite[2][65][29] = 1;dino_sprite[2][65][30] = 1;dino_sprite[2][65][31] = 1;dino_sprite[2][65][32] = 1;dino_sprite[2][65][33] = 1;dino_sprite[2][65][34] = 1;dino_sprite[2][65][35] = 1;dino_sprite[2][65][36] = 1;dino_sprite[2][65][37] = 1;dino_sprite[2][65][38] = 1;dino_sprite[2][65][39] = 1;dino_sprite[2][65][40] = 1;dino_sprite[2][65][41] = 1;dino_sprite[2][65][42] = 1;dino_sprite[2][65][43] = 1;dino_sprite[2][65][44] = 1;dino_sprite[2][65][45] = 1;dino_sprite[2][65][46] = 1;dino_sprite[2][65][47] = 1;dino_sprite[2][65][48] = 1;dino_sprite[2][65][49] = 1;dino_sprite[2][65][50] = 1;dino_sprite[2][65][51] = 1;dino_sprite[2][65][52] = 1;dino_sprite[2][65][53] = 1;dino_sprite[2][65][54] = 1;dino_sprite[2][65][55] = 1;dino_sprite[2][65][56] = 1;dino_sprite[2][65][57] = 1;dino_sprite[2][65][58] = 1;dino_sprite[2][65][59] = 1;dino_sprite[2][65][60] = 1;dino_sprite[2][65][61] = 1;dino_sprite[2][65][62] = 1;dino_sprite[2][65][63] = 1;dino_sprite[2][65][64] = 1;dino_sprite[2][65][65] = 1;dino_sprite[2][65][66] = 1;dino_sprite[2][65][67] = 1;dino_sprite[2][65][68] = 1;dino_sprite[2][65][69] = 1;dino_sprite[2][65][70] = 1;dino_sprite[2][65][71] = 1;dino_sprite[2][65][72] = 1;dino_sprite[2][66][0] = 1;dino_sprite[2][66][1] = 1;dino_sprite[2][66][2] = 1;dino_sprite[2][66][3] = 1;dino_sprite[2][66][4] = 1;dino_sprite[2][66][5] = 1;dino_sprite[2][66][6] = 1;dino_sprite[2][66][7] = 1;dino_sprite[2][66][8] = 1;dino_sprite[2][66][9] = 1;dino_sprite[2][66][10] = 1;dino_sprite[2][66][11] = 1;dino_sprite[2][66][12] = 1;dino_sprite[2][66][13] = 1;dino_sprite[2][66][14] = 1;dino_sprite[2][66][15] = 1;dino_sprite[2][66][16] = 1;dino_sprite[2][66][17] = 1;dino_sprite[2][66][18] = 1;dino_sprite[2][66][19] = 1;dino_sprite[2][66][20] = 1;dino_sprite[2][66][21] = 1;dino_sprite[2][66][22] = 1;dino_sprite[2][66][23] = 1;dino_sprite[2][66][24] = 1;dino_sprite[2][66][25] = 1;dino_sprite[2][66][26] = 1;dino_sprite[2][66][27] = 1;dino_sprite[2][66][28] = 1;dino_sprite[2][66][29] = 1;dino_sprite[2][66][30] = 1;dino_sprite[2][66][31] = 1;dino_sprite[2][66][32] = 1;dino_sprite[2][66][33] = 1;dino_sprite[2][66][34] = 1;dino_sprite[2][66][35] = 1;dino_sprite[2][66][36] = 1;dino_sprite[2][66][37] = 1;dino_sprite[2][66][38] = 1;dino_sprite[2][66][39] = 1;dino_sprite[2][66][40] = 1;dino_sprite[2][66][41] = 1;dino_sprite[2][66][42] = 1;dino_sprite[2][66][43] = 1;dino_sprite[2][66][44] = 1;dino_sprite[2][66][45] = 1;dino_sprite[2][66][46] = 1;dino_sprite[2][66][47] = 1;dino_sprite[2][66][48] = 1;dino_sprite[2][66][49] = 1;dino_sprite[2][66][50] = 1;dino_sprite[2][66][51] = 1;dino_sprite[2][66][52] = 1;dino_sprite[2][66][53] = 1;dino_sprite[2][66][54] = 1;dino_sprite[2][66][55] = 1;dino_sprite[2][66][56] = 1;dino_sprite[2][66][57] = 1;dino_sprite[2][66][58] = 1;dino_sprite[2][66][59] = 1;dino_sprite[2][66][60] = 1;dino_sprite[2][66][61] = 1;dino_sprite[2][66][62] = 1;dino_sprite[2][66][63] = 1;dino_sprite[2][66][64] = 1;dino_sprite[2][66][65] = 1;dino_sprite[2][67][0] = 1;dino_sprite[2][67][1] = 1;dino_sprite[2][67][2] = 1;dino_sprite[2][67][3] = 1;dino_sprite[2][67][4] = 1;dino_sprite[2][67][5] = 1;dino_sprite[2][67][6] = 1;dino_sprite[2][67][7] = 1;dino_sprite[2][67][8] = 1;dino_sprite[2][67][9] = 1;dino_sprite[2][67][10] = 1;dino_sprite[2][67][11] = 1;dino_sprite[2][67][12] = 1;dino_sprite[2][67][13] = 1;dino_sprite[2][67][14] = 1;dino_sprite[2][67][15] = 1;dino_sprite[2][67][16] = 1;dino_sprite[2][67][17] = 1;dino_sprite[2][67][18] = 1;dino_sprite[2][67][19] = 1;dino_sprite[2][67][20] = 1;dino_sprite[2][67][21] = 1;dino_sprite[2][67][22] = 1;dino_sprite[2][67][23] = 1;dino_sprite[2][67][24] = 1;dino_sprite[2][67][25] = 1;dino_sprite[2][67][26] = 1;dino_sprite[2][67][27] = 1;dino_sprite[2][67][28] = 1;dino_sprite[2][67][29] = 1;dino_sprite[2][67][30] = 1;dino_sprite[2][67][31] = 1;dino_sprite[2][67][32] = 1;dino_sprite[2][67][33] = 1;dino_sprite[2][67][34] = 1;dino_sprite[2][67][35] = 1;dino_sprite[2][67][36] = 1;dino_sprite[2][67][37] = 1;dino_sprite[2][67][38] = 1;dino_sprite[2][67][39] = 1;dino_sprite[2][67][40] = 1;dino_sprite[2][67][41] = 1;dino_sprite[2][67][42] = 1;dino_sprite[2][67][43] = 1;dino_sprite[2][67][44] = 1;dino_sprite[2][67][45] = 1;dino_sprite[2][67][46] = 1;dino_sprite[2][67][47] = 1;dino_sprite[2][67][48] = 1;dino_sprite[2][67][49] = 1;dino_sprite[2][67][50] = 1;dino_sprite[2][67][51] = 1;dino_sprite[2][67][52] = 1;dino_sprite[2][67][53] = 1;dino_sprite[2][67][54] = 1;dino_sprite[2][67][55] = 1;dino_sprite[2][67][56] = 1;dino_sprite[2][67][57] = 1;dino_sprite[2][67][58] = 1;dino_sprite[2][67][59] = 1;dino_sprite[2][67][60] = 1;dino_sprite[2][67][61] = 1;dino_sprite[2][67][62] = 1;dino_sprite[2][67][63] = 1;dino_sprite[2][67][64] = 1;dino_sprite[2][67][65] = 1;dino_sprite[2][68][0] = 1;dino_sprite[2][68][1] = 1;dino_sprite[2][68][2] = 1;dino_sprite[2][68][3] = 1;dino_sprite[2][68][4] = 1;dino_sprite[2][68][5] = 1;dino_sprite[2][68][6] = 1;dino_sprite[2][68][7] = 1;dino_sprite[2][68][8] = 1;dino_sprite[2][68][9] = 1;dino_sprite[2][68][10] = 1;dino_sprite[2][68][11] = 1;dino_sprite[2][68][12] = 1;dino_sprite[2][68][13] = 1;dino_sprite[2][68][14] = 1;dino_sprite[2][68][15] = 1;dino_sprite[2][68][16] = 1;dino_sprite[2][68][17] = 1;dino_sprite[2][68][18] = 1;dino_sprite[2][68][19] = 1;dino_sprite[2][68][20] = 1;dino_sprite[2][68][21] = 1;dino_sprite[2][68][22] = 1;dino_sprite[2][68][23] = 1;dino_sprite[2][68][24] = 1;dino_sprite[2][68][25] = 1;dino_sprite[2][68][26] = 1;dino_sprite[2][68][27] = 1;dino_sprite[2][68][28] = 1;dino_sprite[2][68][29] = 1;dino_sprite[2][68][30] = 1;dino_sprite[2][68][31] = 1;dino_sprite[2][68][32] = 1;dino_sprite[2][68][33] = 1;dino_sprite[2][68][34] = 1;dino_sprite[2][68][35] = 1;dino_sprite[2][68][36] = 1;dino_sprite[2][68][37] = 1;dino_sprite[2][68][38] = 1;dino_sprite[2][68][39] = 1;dino_sprite[2][68][40] = 1;dino_sprite[2][68][41] = 1;dino_sprite[2][68][42] = 1;dino_sprite[2][68][43] = 1;dino_sprite[2][68][44] = 1;dino_sprite[2][68][45] = 1;dino_sprite[2][68][46] = 1;dino_sprite[2][68][47] = 1;dino_sprite[2][68][48] = 1;dino_sprite[2][68][49] = 1;dino_sprite[2][68][50] = 1;dino_sprite[2][68][51] = 1;dino_sprite[2][68][52] = 1;dino_sprite[2][68][53] = 1;dino_sprite[2][68][54] = 1;dino_sprite[2][68][55] = 1;dino_sprite[2][68][56] = 1;dino_sprite[2][68][57] = 1;dino_sprite[2][68][58] = 1;dino_sprite[2][68][59] = 1;dino_sprite[2][68][60] = 1;dino_sprite[2][68][61] = 1;dino_sprite[2][68][62] = 1;dino_sprite[2][68][63] = 1;dino_sprite[2][68][64] = 1;dino_sprite[2][68][65] = 1;dino_sprite[2][69][0] = 1;dino_sprite[2][69][1] = 1;dino_sprite[2][69][2] = 1;dino_sprite[2][69][3] = 1;dino_sprite[2][69][4] = 1;dino_sprite[2][69][5] = 1;dino_sprite[2][69][6] = 1;dino_sprite[2][69][7] = 1;dino_sprite[2][69][8] = 1;dino_sprite[2][69][9] = 1;dino_sprite[2][69][10] = 1;dino_sprite[2][69][11] = 1;dino_sprite[2][69][12] = 1;dino_sprite[2][69][13] = 1;dino_sprite[2][69][14] = 1;dino_sprite[2][69][15] = 1;dino_sprite[2][69][16] = 1;dino_sprite[2][69][17] = 1;dino_sprite[2][69][18] = 1;dino_sprite[2][69][19] = 1;dino_sprite[2][69][20] = 1;dino_sprite[2][69][21] = 1;dino_sprite[2][69][22] = 1;dino_sprite[2][69][23] = 1;dino_sprite[2][69][24] = 1;dino_sprite[2][69][25] = 1;dino_sprite[2][69][26] = 1;dino_sprite[2][69][27] = 1;dino_sprite[2][69][28] = 1;dino_sprite[2][69][29] = 1;dino_sprite[2][69][30] = 1;dino_sprite[2][69][31] = 1;dino_sprite[2][69][32] = 1;dino_sprite[2][69][33] = 1;dino_sprite[2][69][34] = 1;dino_sprite[2][69][35] = 1;dino_sprite[2][69][36] = 1;dino_sprite[2][69][37] = 1;dino_sprite[2][69][38] = 1;dino_sprite[2][69][39] = 1;dino_sprite[2][69][40] = 1;dino_sprite[2][69][41] = 1;dino_sprite[2][69][42] = 1;dino_sprite[2][69][43] = 1;dino_sprite[2][69][44] = 1;dino_sprite[2][69][45] = 1;dino_sprite[2][69][46] = 1;dino_sprite[2][69][47] = 1;dino_sprite[2][69][48] = 1;dino_sprite[2][69][49] = 1;dino_sprite[2][69][50] = 1;dino_sprite[2][69][51] = 1;dino_sprite[2][69][52] = 1;dino_sprite[2][69][53] = 1;dino_sprite[2][69][54] = 1;dino_sprite[2][69][55] = 1;dino_sprite[2][69][56] = 1;dino_sprite[2][69][57] = 1;dino_sprite[2][69][58] = 1;dino_sprite[2][69][59] = 1;dino_sprite[2][69][60] = 1;dino_sprite[2][69][61] = 1;dino_sprite[2][69][62] = 1;dino_sprite[2][69][63] = 1;dino_sprite[2][69][64] = 1;dino_sprite[2][69][65] = 1;dino_sprite[2][70][0] = 1;dino_sprite[2][70][1] = 1;dino_sprite[2][70][2] = 1;dino_sprite[2][70][3] = 1;dino_sprite[2][70][4] = 1;dino_sprite[2][70][5] = 1;dino_sprite[2][70][6] = 1;dino_sprite[2][70][7] = 1;dino_sprite[2][70][8] = 1;dino_sprite[2][70][9] = 1;dino_sprite[2][70][10] = 1;dino_sprite[2][70][11] = 1;dino_sprite[2][70][12] = 1;dino_sprite[2][70][13] = 1;dino_sprite[2][70][14] = 1;dino_sprite[2][70][15] = 1;dino_sprite[2][70][16] = 1;dino_sprite[2][70][17] = 1;dino_sprite[2][70][18] = 1;dino_sprite[2][70][19] = 1;dino_sprite[2][70][20] = 1;dino_sprite[2][70][21] = 1;dino_sprite[2][70][22] = 1;dino_sprite[2][70][23] = 1;dino_sprite[2][70][24] = 1;dino_sprite[2][70][25] = 1;dino_sprite[2][70][26] = 1;dino_sprite[2][70][27] = 1;dino_sprite[2][70][28] = 1;dino_sprite[2][70][29] = 1;dino_sprite[2][70][30] = 1;dino_sprite[2][70][31] = 1;dino_sprite[2][70][32] = 1;dino_sprite[2][70][33] = 1;dino_sprite[2][70][34] = 1;dino_sprite[2][70][35] = 1;dino_sprite[2][70][36] = 1;dino_sprite[2][70][37] = 1;dino_sprite[2][70][38] = 1;dino_sprite[2][70][39] = 1;dino_sprite[2][70][40] = 1;dino_sprite[2][70][41] = 1;dino_sprite[2][70][42] = 1;dino_sprite[2][70][43] = 1;dino_sprite[2][70][44] = 1;dino_sprite[2][70][45] = 1;dino_sprite[2][70][46] = 1;dino_sprite[2][70][47] = 1;dino_sprite[2][70][48] = 1;dino_sprite[2][70][49] = 1;dino_sprite[2][70][50] = 1;dino_sprite[2][70][51] = 1;dino_sprite[2][70][52] = 1;dino_sprite[2][70][53] = 1;dino_sprite[2][70][54] = 1;dino_sprite[2][70][55] = 1;dino_sprite[2][70][56] = 1;dino_sprite[2][70][57] = 1;dino_sprite[2][70][58] = 1;dino_sprite[2][70][59] = 1;dino_sprite[2][70][60] = 1;dino_sprite[2][70][61] = 1;dino_sprite[2][70][62] = 1;dino_sprite[2][70][63] = 1;dino_sprite[2][70][64] = 1;dino_sprite[2][70][65] = 1;dino_sprite[2][71][0] = 1;dino_sprite[2][71][1] = 1;dino_sprite[2][71][2] = 1;dino_sprite[2][71][3] = 1;dino_sprite[2][71][4] = 1;dino_sprite[2][71][5] = 1;dino_sprite[2][71][6] = 1;dino_sprite[2][71][7] = 1;dino_sprite[2][71][8] = 1;dino_sprite[2][71][9] = 1;dino_sprite[2][71][10] = 1;dino_sprite[2][71][11] = 1;dino_sprite[2][71][12] = 1;dino_sprite[2][71][13] = 1;dino_sprite[2][71][14] = 1;dino_sprite[2][71][15] = 1;dino_sprite[2][71][16] = 1;dino_sprite[2][71][17] = 1;dino_sprite[2][71][18] = 1;dino_sprite[2][71][19] = 1;dino_sprite[2][71][20] = 1;dino_sprite[2][71][21] = 1;dino_sprite[2][71][22] = 1;dino_sprite[2][71][23] = 1;dino_sprite[2][71][24] = 1;dino_sprite[2][71][25] = 1;dino_sprite[2][71][26] = 1;dino_sprite[2][71][27] = 1;dino_sprite[2][71][28] = 1;dino_sprite[2][71][29] = 1;dino_sprite[2][71][30] = 1;dino_sprite[2][71][31] = 1;dino_sprite[2][71][32] = 1;dino_sprite[2][71][33] = 1;dino_sprite[2][71][34] = 1;dino_sprite[2][71][35] = 1;dino_sprite[2][71][36] = 1;dino_sprite[2][71][37] = 1;dino_sprite[2][71][38] = 1;dino_sprite[2][71][39] = 1;dino_sprite[2][71][40] = 1;dino_sprite[2][71][41] = 1;dino_sprite[2][71][43] = 1;dino_sprite[2][71][44] = 1;dino_sprite[2][71][45] = 1;dino_sprite[2][71][46] = 1;dino_sprite[2][71][47] = 1;dino_sprite[2][71][48] = 1;dino_sprite[2][71][49] = 1;dino_sprite[2][72][0] = 1;dino_sprite[2][72][1] = 1;dino_sprite[2][72][2] = 1;dino_sprite[2][72][3] = 1;dino_sprite[2][72][4] = 1;dino_sprite[2][72][5] = 1;dino_sprite[2][72][6] = 1;dino_sprite[2][72][7] = 1;dino_sprite[2][72][8] = 1;dino_sprite[2][72][9] = 1;dino_sprite[2][72][10] = 1;dino_sprite[2][72][11] = 1;dino_sprite[2][72][12] = 1;dino_sprite[2][72][13] = 1;dino_sprite[2][72][14] = 1;dino_sprite[2][72][15] = 1;dino_sprite[2][72][16] = 1;dino_sprite[2][72][17] = 1;dino_sprite[2][72][18] = 1;dino_sprite[2][72][19] = 1;dino_sprite[2][72][20] = 1;dino_sprite[2][72][21] = 1;dino_sprite[2][72][22] = 1;dino_sprite[2][72][23] = 1;dino_sprite[2][72][24] = 1;dino_sprite[2][72][25] = 1;dino_sprite[2][72][26] = 1;dino_sprite[2][72][27] = 1;dino_sprite[2][72][28] = 1;dino_sprite[2][72][29] = 1;dino_sprite[2][72][30] = 1;dino_sprite[2][72][31] = 1;dino_sprite[2][72][32] = 1;dino_sprite[2][72][33] = 1;dino_sprite[2][72][34] = 1;dino_sprite[2][72][35] = 1;dino_sprite[2][72][43] = 1;dino_sprite[2][72][44] = 1;dino_sprite[2][72][45] = 1;dino_sprite[2][72][46] = 1;dino_sprite[2][72][47] = 1;dino_sprite[2][72][48] = 1;dino_sprite[2][72][49] = 1;dino_sprite[2][73][0] = 1;dino_sprite[2][73][1] = 1;dino_sprite[2][73][2] = 1;dino_sprite[2][73][3] = 1;dino_sprite[2][73][4] = 1;dino_sprite[2][73][5] = 1;dino_sprite[2][73][6] = 1;dino_sprite[2][73][7] = 1;dino_sprite[2][73][8] = 1;dino_sprite[2][73][9] = 1;dino_sprite[2][73][10] = 1;dino_sprite[2][73][11] = 1;dino_sprite[2][73][12] = 1;dino_sprite[2][73][13] = 1;dino_sprite[2][73][14] = 1;dino_sprite[2][73][15] = 1;dino_sprite[2][73][16] = 1;dino_sprite[2][73][17] = 1;dino_sprite[2][73][18] = 1;dino_sprite[2][73][19] = 1;dino_sprite[2][73][20] = 1;dino_sprite[2][73][21] = 1;dino_sprite[2][73][22] = 1;dino_sprite[2][73][23] = 1;dino_sprite[2][73][24] = 1;dino_sprite[2][73][25] = 1;dino_sprite[2][73][26] = 1;dino_sprite[2][73][27] = 1;dino_sprite[2][73][28] = 1;dino_sprite[2][73][29] = 1;dino_sprite[2][73][30] = 1;dino_sprite[2][73][31] = 1;dino_sprite[2][73][32] = 1;dino_sprite[2][73][33] = 1;dino_sprite[2][73][34] = 1;dino_sprite[2][73][35] = 1;dino_sprite[2][73][43] = 1;dino_sprite[2][73][44] = 1;dino_sprite[2][73][45] = 1;dino_sprite[2][73][46] = 1;dino_sprite[2][73][47] = 1;dino_sprite[2][73][48] = 1;dino_sprite[2][73][49] = 1;dino_sprite[2][74][0] = 1;dino_sprite[2][74][1] = 1;dino_sprite[2][74][2] = 1;dino_sprite[2][74][3] = 1;dino_sprite[2][74][4] = 1;dino_sprite[2][74][5] = 1;dino_sprite[2][74][6] = 1;dino_sprite[2][74][7] = 1;dino_sprite[2][74][8] = 1;dino_sprite[2][74][9] = 1;dino_sprite[2][74][10] = 1;dino_sprite[2][74][11] = 1;dino_sprite[2][74][12] = 1;dino_sprite[2][74][13] = 1;dino_sprite[2][74][14] = 1;dino_sprite[2][74][15] = 1;dino_sprite[2][74][16] = 1;dino_sprite[2][74][17] = 1;dino_sprite[2][74][18] = 1;dino_sprite[2][74][19] = 1;dino_sprite[2][74][20] = 1;dino_sprite[2][74][21] = 1;dino_sprite[2][74][22] = 1;dino_sprite[2][74][23] = 1;dino_sprite[2][74][24] = 1;dino_sprite[2][74][25] = 1;dino_sprite[2][74][26] = 1;dino_sprite[2][74][27] = 1;dino_sprite[2][74][28] = 1;dino_sprite[2][74][29] = 1;dino_sprite[2][74][30] = 1;dino_sprite[2][74][31] = 1;dino_sprite[2][74][32] = 1;dino_sprite[2][74][33] = 1;dino_sprite[2][74][34] = 1;dino_sprite[2][74][35] = 1;dino_sprite[2][74][43] = 1;dino_sprite[2][74][44] = 1;dino_sprite[2][74][45] = 1;dino_sprite[2][74][46] = 1;dino_sprite[2][74][47] = 1;dino_sprite[2][74][48] = 1;dino_sprite[2][74][49] = 1;dino_sprite[2][75][0] = 1;dino_sprite[2][75][1] = 1;dino_sprite[2][75][2] = 1;dino_sprite[2][75][3] = 1;dino_sprite[2][75][4] = 1;dino_sprite[2][75][5] = 1;dino_sprite[2][75][6] = 1;dino_sprite[2][75][7] = 1;dino_sprite[2][75][8] = 1;dino_sprite[2][75][9] = 1;dino_sprite[2][75][10] = 1;dino_sprite[2][75][11] = 1;dino_sprite[2][75][12] = 1;dino_sprite[2][75][13] = 1;dino_sprite[2][75][14] = 1;dino_sprite[2][75][15] = 1;dino_sprite[2][75][16] = 1;dino_sprite[2][75][17] = 1;dino_sprite[2][75][18] = 1;dino_sprite[2][75][19] = 1;dino_sprite[2][75][20] = 1;dino_sprite[2][75][21] = 1;dino_sprite[2][75][22] = 1;dino_sprite[2][75][23] = 1;dino_sprite[2][75][24] = 1;dino_sprite[2][75][25] = 1;dino_sprite[2][75][26] = 1;dino_sprite[2][75][27] = 1;dino_sprite[2][75][28] = 1;dino_sprite[2][75][29] = 1;dino_sprite[2][75][30] = 1;dino_sprite[2][75][31] = 1;dino_sprite[2][75][32] = 1;dino_sprite[2][75][33] = 1;dino_sprite[2][75][34] = 1;dino_sprite[2][75][35] = 1;dino_sprite[2][75][43] = 1;dino_sprite[2][75][44] = 1;dino_sprite[2][75][45] = 1;dino_sprite[2][75][46] = 1;dino_sprite[2][75][47] = 1;dino_sprite[2][75][48] = 1;dino_sprite[2][75][49] = 1;dino_sprite[2][75][50] = 1;dino_sprite[2][75][51] = 1;dino_sprite[2][75][52] = 1;dino_sprite[2][75][53] = 1;dino_sprite[2][75][54] = 1;dino_sprite[2][76][0] = 1;dino_sprite[2][76][1] = 1;dino_sprite[2][76][2] = 1;dino_sprite[2][76][3] = 1;dino_sprite[2][76][4] = 1;dino_sprite[2][76][5] = 1;dino_sprite[2][76][6] = 1;dino_sprite[2][76][7] = 1;dino_sprite[2][76][8] = 1;dino_sprite[2][76][9] = 1;dino_sprite[2][76][10] = 1;dino_sprite[2][76][11] = 1;dino_sprite[2][76][12] = 1;dino_sprite[2][76][13] = 1;dino_sprite[2][76][14] = 1;dino_sprite[2][76][15] = 1;dino_sprite[2][76][16] = 1;dino_sprite[2][76][17] = 1;dino_sprite[2][76][18] = 1;dino_sprite[2][76][19] = 1;dino_sprite[2][76][20] = 1;dino_sprite[2][76][21] = 1;dino_sprite[2][76][22] = 1;dino_sprite[2][76][23] = 1;dino_sprite[2][76][24] = 1;dino_sprite[2][76][25] = 1;dino_sprite[2][76][26] = 1;dino_sprite[2][76][27] = 1;dino_sprite[2][76][28] = 1;dino_sprite[2][76][29] = 1;dino_sprite[2][76][30] = 1;dino_sprite[2][76][31] = 1;dino_sprite[2][76][32] = 1;dino_sprite[2][76][33] = 1;dino_sprite[2][76][34] = 1;dino_sprite[2][76][35] = 1;dino_sprite[2][76][43] = 1;dino_sprite[2][76][44] = 1;dino_sprite[2][76][45] = 1;dino_sprite[2][76][46] = 1;dino_sprite[2][76][47] = 1;dino_sprite[2][76][48] = 1;dino_sprite[2][76][49] = 1;dino_sprite[2][76][50] = 1;dino_sprite[2][76][51] = 1;dino_sprite[2][76][52] = 1;dino_sprite[2][76][53] = 1;dino_sprite[2][76][54] = 1;dino_sprite[2][77][0] = 1;dino_sprite[2][77][1] = 1;dino_sprite[2][77][2] = 1;dino_sprite[2][77][3] = 1;dino_sprite[2][77][4] = 1;dino_sprite[2][77][5] = 1;dino_sprite[2][77][6] = 1;dino_sprite[2][77][7] = 1;dino_sprite[2][77][8] = 1;dino_sprite[2][77][9] = 1;dino_sprite[2][77][10] = 1;dino_sprite[2][77][11] = 1;dino_sprite[2][77][12] = 1;dino_sprite[2][77][13] = 1;dino_sprite[2][77][14] = 1;dino_sprite[2][77][15] = 1;dino_sprite[2][77][16] = 1;dino_sprite[2][77][17] = 1;dino_sprite[2][77][18] = 1;dino_sprite[2][77][19] = 1;dino_sprite[2][77][20] = 1;dino_sprite[2][77][21] = 1;dino_sprite[2][77][22] = 1;dino_sprite[2][77][23] = 1;dino_sprite[2][77][24] = 1;dino_sprite[2][77][25] = 1;dino_sprite[2][77][29] = 1;dino_sprite[2][77][30] = 1;dino_sprite[2][77][31] = 1;dino_sprite[2][77][32] = 1;dino_sprite[2][77][33] = 1;dino_sprite[2][77][34] = 1;dino_sprite[2][77][35] = 1;dino_sprite[2][77][43] = 1;dino_sprite[2][77][44] = 1;dino_sprite[2][77][45] = 1;dino_sprite[2][77][46] = 1;dino_sprite[2][77][47] = 1;dino_sprite[2][77][48] = 1;dino_sprite[2][77][49] = 1;dino_sprite[2][77][50] = 1;dino_sprite[2][77][51] = 1;dino_sprite[2][77][52] = 1;dino_sprite[2][77][53] = 1;dino_sprite[2][77][54] = 1;dino_sprite[2][78][0] = 1;dino_sprite[2][78][1] = 1;dino_sprite[2][78][2] = 1;dino_sprite[2][78][3] = 1;dino_sprite[2][78][4] = 1;dino_sprite[2][78][5] = 1;dino_sprite[2][78][6] = 1;dino_sprite[2][78][7] = 1;dino_sprite[2][78][8] = 1;dino_sprite[2][78][9] = 1;dino_sprite[2][78][10] = 1;dino_sprite[2][78][11] = 1;dino_sprite[2][78][12] = 1;dino_sprite[2][78][13] = 1;dino_sprite[2][78][14] = 1;dino_sprite[2][78][15] = 1;dino_sprite[2][78][16] = 1;dino_sprite[2][78][17] = 1;dino_sprite[2][78][18] = 1;dino_sprite[2][78][19] = 1;dino_sprite[2][78][20] = 1;dino_sprite[2][78][21] = 1;dino_sprite[2][78][22] = 1;dino_sprite[2][78][23] = 1;dino_sprite[2][78][24] = 1;dino_sprite[2][78][25] = 1;dino_sprite[2][78][29] = 1;dino_sprite[2][78][30] = 1;dino_sprite[2][78][31] = 1;dino_sprite[2][78][32] = 1;dino_sprite[2][78][33] = 1;dino_sprite[2][78][34] = 1;dino_sprite[2][78][35] = 1;dino_sprite[2][78][43] = 1;dino_sprite[2][78][44] = 1;dino_sprite[2][78][45] = 1;dino_sprite[2][78][46] = 1;dino_sprite[2][78][47] = 1;dino_sprite[2][78][48] = 1;dino_sprite[2][78][49] = 1;dino_sprite[2][78][50] = 1;dino_sprite[2][78][51] = 1;dino_sprite[2][78][52] = 1;dino_sprite[2][78][53] = 1;dino_sprite[2][78][54] = 1;dino_sprite[2][79][0] = 1;dino_sprite[2][79][1] = 1;dino_sprite[2][79][2] = 1;dino_sprite[2][79][3] = 1;dino_sprite[2][79][4] = 1;dino_sprite[2][79][5] = 1;dino_sprite[2][79][6] = 1;dino_sprite[2][79][7] = 1;dino_sprite[2][79][8] = 1;dino_sprite[2][79][9] = 1;dino_sprite[2][79][10] = 1;dino_sprite[2][79][11] = 1;dino_sprite[2][79][12] = 1;dino_sprite[2][79][13] = 1;dino_sprite[2][79][14] = 1;dino_sprite[2][79][15] = 1;dino_sprite[2][79][16] = 1;dino_sprite[2][79][17] = 1;dino_sprite[2][79][18] = 1;dino_sprite[2][79][19] = 1;dino_sprite[2][79][20] = 1;dino_sprite[2][79][21] = 1;dino_sprite[2][79][22] = 1;dino_sprite[2][79][23] = 1;dino_sprite[2][79][24] = 1;dino_sprite[2][79][25] = 1;dino_sprite[2][79][29] = 1;dino_sprite[2][79][30] = 1;dino_sprite[2][79][31] = 1;dino_sprite[2][79][32] = 1;dino_sprite[2][79][33] = 1;dino_sprite[2][79][34] = 1;dino_sprite[2][79][35] = 1;dino_sprite[2][79][43] = 1;dino_sprite[2][79][44] = 1;dino_sprite[2][79][45] = 1;dino_sprite[2][79][46] = 1;dino_sprite[2][79][47] = 1;dino_sprite[2][79][48] = 1;dino_sprite[2][79][49] = 1;dino_sprite[2][79][50] = 1;dino_sprite[2][79][51] = 1;dino_sprite[2][79][52] = 1;dino_sprite[2][79][53] = 1;dino_sprite[2][79][54] = 1;dino_sprite[2][80][0] = 1;dino_sprite[2][80][1] = 1;dino_sprite[2][80][2] = 1;dino_sprite[2][80][3] = 1;dino_sprite[2][80][4] = 1;dino_sprite[2][80][5] = 1;dino_sprite[2][80][6] = 1;dino_sprite[2][80][7] = 1;dino_sprite[2][80][8] = 1;dino_sprite[2][80][9] = 1;dino_sprite[2][80][10] = 1;dino_sprite[2][80][11] = 1;dino_sprite[2][80][12] = 1;dino_sprite[2][80][13] = 1;dino_sprite[2][80][14] = 1;dino_sprite[2][80][15] = 1;dino_sprite[2][80][16] = 1;dino_sprite[2][80][17] = 1;dino_sprite[2][80][18] = 1;dino_sprite[2][80][19] = 1;dino_sprite[2][80][20] = 1;dino_sprite[2][80][21] = 1;dino_sprite[2][80][22] = 1;dino_sprite[2][80][23] = 1;dino_sprite[2][80][24] = 1;dino_sprite[2][80][25] = 1;dino_sprite[2][80][29] = 1;dino_sprite[2][80][30] = 1;dino_sprite[2][80][31] = 1;dino_sprite[2][80][32] = 1;dino_sprite[2][80][33] = 1;dino_sprite[2][80][34] = 1;dino_sprite[2][80][35] = 1;dino_sprite[2][80][43] = 1;dino_sprite[2][80][44] = 1;dino_sprite[2][80][45] = 1;dino_sprite[2][80][46] = 1;dino_sprite[2][80][47] = 1;dino_sprite[2][80][48] = 1;dino_sprite[2][80][49] = 1;dino_sprite[2][80][50] = 1;dino_sprite[2][80][51] = 1;dino_sprite[2][80][52] = 1;dino_sprite[2][80][53] = 1;dino_sprite[2][80][54] = 1;dino_sprite[2][81][0] = 1;dino_sprite[2][81][1] = 1;dino_sprite[2][81][2] = 1;dino_sprite[2][81][3] = 1;dino_sprite[2][81][4] = 1;dino_sprite[2][81][5] = 1;dino_sprite[2][81][6] = 1;dino_sprite[2][81][7] = 1;dino_sprite[2][81][8] = 1;dino_sprite[2][81][9] = 1;dino_sprite[2][81][10] = 1;dino_sprite[2][81][11] = 1;dino_sprite[2][81][12] = 1;dino_sprite[2][81][13] = 1;dino_sprite[2][81][14] = 1;dino_sprite[2][81][15] = 1;dino_sprite[2][81][16] = 1;dino_sprite[2][81][17] = 1;dino_sprite[2][81][18] = 1;dino_sprite[2][81][19] = 1;dino_sprite[2][81][20] = 1;dino_sprite[2][81][21] = 1;dino_sprite[2][81][22] = 1;dino_sprite[2][81][23] = 1;dino_sprite[2][81][24] = 1;dino_sprite[2][81][25] = 1;dino_sprite[2][81][29] = 1;dino_sprite[2][81][30] = 1;dino_sprite[2][81][31] = 1;dino_sprite[2][81][32] = 1;dino_sprite[2][81][33] = 1;dino_sprite[2][81][34] = 1;dino_sprite[2][81][35] = 1;dino_sprite[2][81][43] = 1;dino_sprite[2][81][44] = 1;dino_sprite[2][81][45] = 1;dino_sprite[2][81][46] = 1;dino_sprite[2][81][47] = 1;dino_sprite[2][81][48] = 1;dino_sprite[2][81][49] = 1;dino_sprite[2][81][50] = 1;dino_sprite[2][81][51] = 1;dino_sprite[2][81][52] = 1;dino_sprite[2][81][53] = 1;dino_sprite[2][81][54] = 1;dino_sprite[2][82][0] = 1;dino_sprite[2][82][1] = 1;dino_sprite[2][82][2] = 1;dino_sprite[2][82][3] = 1;dino_sprite[2][82][4] = 1;dino_sprite[2][82][5] = 1;dino_sprite[2][82][6] = 1;dino_sprite[2][82][7] = 1;dino_sprite[2][82][8] = 1;dino_sprite[2][82][9] = 1;dino_sprite[2][82][10] = 1;dino_sprite[2][82][11] = 1;dino_sprite[2][82][12] = 1;dino_sprite[2][82][13] = 1;dino_sprite[2][82][14] = 1;dino_sprite[2][82][15] = 1;dino_sprite[2][82][16] = 1;dino_sprite[2][82][17] = 1;dino_sprite[2][82][18] = 1;dino_sprite[2][82][19] = 1;dino_sprite[2][82][20] = 1;dino_sprite[2][82][21] = 1;dino_sprite[2][82][22] = 1;dino_sprite[2][82][23] = 1;dino_sprite[2][82][24] = 1;dino_sprite[2][82][25] = 1;dino_sprite[2][82][29] = 1;dino_sprite[2][82][30] = 1;dino_sprite[2][82][31] = 1;dino_sprite[2][82][32] = 1;dino_sprite[2][82][33] = 1;dino_sprite[2][82][34] = 1;dino_sprite[2][82][35] = 1;dino_sprite[2][83][0] = 1;dino_sprite[2][83][1] = 1;dino_sprite[2][83][2] = 1;dino_sprite[2][83][3] = 1;dino_sprite[2][83][4] = 1;dino_sprite[2][83][5] = 1;dino_sprite[2][83][6] = 1;dino_sprite[2][83][7] = 1;dino_sprite[2][83][8] = 1;dino_sprite[2][83][9] = 1;dino_sprite[2][83][10] = 1;dino_sprite[2][83][11] = 1;dino_sprite[2][83][12] = 1;dino_sprite[2][83][13] = 1;dino_sprite[2][83][14] = 1;dino_sprite[2][83][15] = 1;dino_sprite[2][83][16] = 1;dino_sprite[2][83][17] = 1;dino_sprite[2][83][18] = 1;dino_sprite[2][83][19] = 1;dino_sprite[2][83][20] = 1;dino_sprite[2][83][21] = 1;dino_sprite[2][83][22] = 1;dino_sprite[2][83][23] = 1;dino_sprite[2][83][24] = 1;dino_sprite[2][83][25] = 1;dino_sprite[2][83][29] = 1;dino_sprite[2][83][30] = 1;dino_sprite[2][83][31] = 1;dino_sprite[2][83][32] = 1;dino_sprite[2][83][33] = 1;dino_sprite[2][83][34] = 1;dino_sprite[2][83][35] = 1;dino_sprite[2][84][0] = 1;dino_sprite[2][84][1] = 1;dino_sprite[2][84][2] = 1;dino_sprite[2][84][3] = 1;dino_sprite[2][84][4] = 1;dino_sprite[2][84][5] = 1;dino_sprite[2][84][6] = 1;dino_sprite[2][84][7] = 1;dino_sprite[2][84][8] = 1;dino_sprite[2][84][9] = 1;dino_sprite[2][84][10] = 1;dino_sprite[2][84][11] = 1;dino_sprite[2][84][12] = 1;dino_sprite[2][84][13] = 1;dino_sprite[2][84][14] = 1;dino_sprite[2][84][15] = 1;dino_sprite[2][84][16] = 1;dino_sprite[2][84][17] = 1;dino_sprite[2][84][18] = 1;dino_sprite[2][84][19] = 1;dino_sprite[2][84][20] = 1;dino_sprite[2][84][21] = 1;dino_sprite[2][84][22] = 1;dino_sprite[2][84][23] = 1;dino_sprite[2][84][24] = 1;dino_sprite[2][84][25] = 1;dino_sprite[2][84][29] = 1;dino_sprite[2][84][30] = 1;dino_sprite[2][84][31] = 1;dino_sprite[2][84][32] = 1;dino_sprite[2][84][33] = 1;dino_sprite[2][84][34] = 1;dino_sprite[2][84][35] = 1;dino_sprite[2][85][0] = 1;dino_sprite[2][85][1] = 1;dino_sprite[2][85][2] = 1;dino_sprite[2][85][3] = 1;dino_sprite[2][85][4] = 1;dino_sprite[2][85][5] = 1;dino_sprite[2][85][6] = 1;dino_sprite[2][85][7] = 1;dino_sprite[2][85][8] = 1;dino_sprite[2][85][9] = 1;dino_sprite[2][85][10] = 1;dino_sprite[2][85][11] = 1;dino_sprite[2][85][12] = 1;dino_sprite[2][85][13] = 1;dino_sprite[2][85][14] = 1;dino_sprite[2][85][15] = 1;dino_sprite[2][85][16] = 1;dino_sprite[2][85][17] = 1;dino_sprite[2][85][18] = 1;dino_sprite[2][85][19] = 1;dino_sprite[2][85][20] = 1;dino_sprite[2][85][21] = 1;dino_sprite[2][85][22] = 1;dino_sprite[2][85][23] = 1;dino_sprite[2][85][24] = 1;dino_sprite[2][85][25] = 1;dino_sprite[2][85][29] = 1;dino_sprite[2][85][30] = 1;dino_sprite[2][85][31] = 1;dino_sprite[2][85][32] = 1;dino_sprite[2][85][33] = 1;dino_sprite[2][85][34] = 1;dino_sprite[2][85][35] = 1;dino_sprite[2][86][0] = 1;dino_sprite[2][86][1] = 1;dino_sprite[2][86][2] = 1;dino_sprite[2][86][3] = 1;dino_sprite[2][86][4] = 1;dino_sprite[2][86][5] = 1;dino_sprite[2][86][6] = 1;dino_sprite[2][86][7] = 1;dino_sprite[2][86][8] = 1;dino_sprite[2][86][9] = 1;dino_sprite[2][86][10] = 1;dino_sprite[2][86][11] = 1;dino_sprite[2][86][12] = 1;dino_sprite[2][86][13] = 1;dino_sprite[2][86][14] = 1;dino_sprite[2][86][15] = 1;dino_sprite[2][86][16] = 1;dino_sprite[2][86][17] = 1;dino_sprite[2][86][18] = 1;dino_sprite[2][86][19] = 1;dino_sprite[2][86][20] = 1;dino_sprite[2][86][21] = 1;dino_sprite[2][86][22] = 1;dino_sprite[2][86][23] = 1;dino_sprite[2][86][24] = 1;dino_sprite[2][86][25] = 1;dino_sprite[2][86][29] = 1;dino_sprite[2][86][30] = 1;dino_sprite[2][86][31] = 1;dino_sprite[2][86][32] = 1;dino_sprite[2][86][33] = 1;dino_sprite[2][86][34] = 1;dino_sprite[2][86][35] = 1;dino_sprite[2][87][0] = 1;dino_sprite[2][87][1] = 1;dino_sprite[2][87][2] = 1;dino_sprite[2][87][3] = 1;dino_sprite[2][87][4] = 1;dino_sprite[2][87][5] = 1;dino_sprite[2][87][6] = 1;dino_sprite[2][87][7] = 1;dino_sprite[2][87][8] = 1;dino_sprite[2][87][9] = 1;dino_sprite[2][87][10] = 1;dino_sprite[2][87][11] = 1;dino_sprite[2][87][12] = 1;dino_sprite[2][87][13] = 1;dino_sprite[2][87][14] = 1;dino_sprite[2][87][15] = 1;dino_sprite[2][87][16] = 1;dino_sprite[2][87][17] = 1;dino_sprite[2][87][18] = 1;dino_sprite[2][87][19] = 1;dino_sprite[2][87][20] = 1;dino_sprite[2][87][21] = 1;dino_sprite[2][87][22] = 1;dino_sprite[2][87][23] = 1;dino_sprite[2][87][24] = 1;dino_sprite[2][87][25] = 1;dino_sprite[2][87][29] = 1;dino_sprite[2][87][30] = 1;dino_sprite[2][87][31] = 1;dino_sprite[2][87][32] = 1;dino_sprite[2][87][33] = 1;dino_sprite[2][87][34] = 1;dino_sprite[2][87][35] = 1;dino_sprite[2][88][0] = 1;dino_sprite[2][88][1] = 1;dino_sprite[2][88][2] = 1;dino_sprite[2][88][3] = 1;dino_sprite[2][88][4] = 1;dino_sprite[2][88][5] = 1;dino_sprite[2][88][6] = 1;dino_sprite[2][88][7] = 1;dino_sprite[2][88][8] = 1;dino_sprite[2][88][9] = 1;dino_sprite[2][88][10] = 1;dino_sprite[2][88][11] = 1;dino_sprite[2][88][12] = 1;dino_sprite[2][88][13] = 1;dino_sprite[2][88][14] = 1;dino_sprite[2][88][15] = 1;dino_sprite[2][88][16] = 1;dino_sprite[2][88][17] = 1;dino_sprite[2][88][18] = 1;dino_sprite[2][88][19] = 1;dino_sprite[2][88][20] = 1;dino_sprite[2][88][21] = 1;dino_sprite[2][88][22] = 1;dino_sprite[2][88][23] = 1;dino_sprite[2][88][24] = 1;dino_sprite[2][88][25] = 1;dino_sprite[2][88][29] = 1;dino_sprite[2][88][30] = 1;dino_sprite[2][88][31] = 1;dino_sprite[2][88][32] = 1;dino_sprite[2][88][33] = 1;dino_sprite[2][88][34] = 1;dino_sprite[2][88][35] = 1;dino_sprite[2][89][0] = 1;dino_sprite[2][89][1] = 1;dino_sprite[2][89][2] = 1;dino_sprite[2][89][3] = 1;dino_sprite[2][89][4] = 1;dino_sprite[2][89][5] = 1;dino_sprite[2][89][6] = 1;dino_sprite[2][89][7] = 1;dino_sprite[2][89][8] = 1;dino_sprite[2][89][9] = 1;dino_sprite[2][89][10] = 1;dino_sprite[2][89][11] = 1;dino_sprite[2][89][12] = 1;dino_sprite[2][89][13] = 1;dino_sprite[2][89][14] = 1;dino_sprite[2][89][15] = 1;dino_sprite[2][89][16] = 1;dino_sprite[2][89][17] = 1;dino_sprite[2][89][18] = 1;dino_sprite[2][89][19] = 1;dino_sprite[2][89][20] = 1;dino_sprite[2][89][21] = 1;dino_sprite[2][89][22] = 1;dino_sprite[2][89][23] = 1;dino_sprite[2][89][24] = 1;dino_sprite[2][89][25] = 1;dino_sprite[2][89][29] = 1;dino_sprite[2][89][30] = 1;dino_sprite[2][89][31] = 1;dino_sprite[2][89][32] = 1;dino_sprite[2][89][33] = 1;dino_sprite[2][89][34] = 1;dino_sprite[2][89][35] = 1;dino_sprite[2][90][0] = 1;dino_sprite[2][90][1] = 1;dino_sprite[2][90][2] = 1;dino_sprite[2][90][3] = 1;dino_sprite[2][90][4] = 1;dino_sprite[2][90][5] = 1;dino_sprite[2][90][6] = 1;dino_sprite[2][90][7] = 1;dino_sprite[2][90][8] = 1;dino_sprite[2][90][9] = 1;dino_sprite[2][90][10] = 1;dino_sprite[2][90][11] = 1;dino_sprite[2][90][12] = 1;dino_sprite[2][90][13] = 1;dino_sprite[2][90][14] = 1;dino_sprite[2][90][15] = 1;dino_sprite[2][90][16] = 1;dino_sprite[2][90][17] = 1;dino_sprite[2][90][18] = 1;dino_sprite[2][90][19] = 1;dino_sprite[2][90][20] = 1;dino_sprite[2][90][21] = 1;dino_sprite[2][90][22] = 1;dino_sprite[2][90][23] = 1;dino_sprite[2][90][24] = 1;dino_sprite[2][90][25] = 1;dino_sprite[2][90][29] = 1;dino_sprite[2][90][30] = 1;dino_sprite[2][90][31] = 1;dino_sprite[2][90][32] = 1;dino_sprite[2][90][33] = 1;dino_sprite[2][90][34] = 1;dino_sprite[2][90][35] = 1;dino_sprite[2][91][0] = 1;dino_sprite[2][91][1] = 1;dino_sprite[2][91][2] = 1;dino_sprite[2][91][3] = 1;dino_sprite[2][91][4] = 1;dino_sprite[2][91][5] = 1;dino_sprite[2][91][6] = 1;dino_sprite[2][91][7] = 1;dino_sprite[2][91][8] = 1;dino_sprite[2][91][9] = 1;dino_sprite[2][91][10] = 1;dino_sprite[2][91][11] = 1;dino_sprite[2][91][12] = 1;dino_sprite[2][91][13] = 1;dino_sprite[2][91][14] = 1;dino_sprite[2][91][15] = 1;dino_sprite[2][91][16] = 1;dino_sprite[2][91][17] = 1;dino_sprite[2][91][18] = 1;dino_sprite[2][91][19] = 1;dino_sprite[2][91][20] = 1;dino_sprite[2][91][21] = 1;dino_sprite[2][91][22] = 1;dino_sprite[2][91][23] = 1;dino_sprite[2][91][24] = 1;dino_sprite[2][91][25] = 1;dino_sprite[2][91][30] = 1;dino_sprite[2][91][31] = 1;dino_sprite[2][91][32] = 1;dino_sprite[2][91][33] = 1;dino_sprite[2][92][0] = 1;dino_sprite[2][92][1] = 1;dino_sprite[2][92][2] = 1;dino_sprite[2][92][3] = 1;dino_sprite[2][92][4] = 1;dino_sprite[2][92][5] = 1;dino_sprite[2][92][6] = 1;dino_sprite[2][92][7] = 1;dino_sprite[2][92][8] = 1;dino_sprite[2][92][9] = 1;dino_sprite[2][92][10] = 1;dino_sprite[2][92][11] = 1;dino_sprite[2][92][12] = 1;dino_sprite[2][92][13] = 1;dino_sprite[2][92][14] = 1;dino_sprite[2][92][15] = 1;dino_sprite[2][92][16] = 1;dino_sprite[2][92][17] = 1;dino_sprite[2][92][18] = 1;dino_sprite[2][92][19] = 1;dino_sprite[2][92][20] = 1;dino_sprite[2][92][21] = 1;dino_sprite[2][92][22] = 1;dino_sprite[2][92][23] = 1;dino_sprite[2][92][24] = 1;dino_sprite[2][92][25] = 1;dino_sprite[2][93][0] = 1;dino_sprite[2][93][1] = 1;dino_sprite[2][93][2] = 1;dino_sprite[2][93][3] = 1;dino_sprite[2][93][4] = 1;dino_sprite[2][93][5] = 1;dino_sprite[2][93][6] = 1;dino_sprite[2][93][7] = 1;dino_sprite[2][93][8] = 1;dino_sprite[2][93][9] = 1;dino_sprite[2][93][10] = 1;dino_sprite[2][93][11] = 1;dino_sprite[2][93][12] = 1;dino_sprite[2][93][13] = 1;dino_sprite[2][93][14] = 1;dino_sprite[2][93][15] = 1;dino_sprite[2][93][16] = 1;dino_sprite[2][93][17] = 1;dino_sprite[2][93][18] = 1;dino_sprite[2][93][19] = 1;dino_sprite[2][93][20] = 1;dino_sprite[2][93][21] = 1;dino_sprite[2][93][22] = 1;dino_sprite[2][93][23] = 1;dino_sprite[2][93][24] = 1;dino_sprite[2][93][25] = 1;dino_sprite[2][94][0] = 1;dino_sprite[2][94][1] = 1;dino_sprite[2][94][2] = 1;dino_sprite[2][94][3] = 1;dino_sprite[2][94][4] = 1;dino_sprite[2][94][5] = 1;dino_sprite[2][94][6] = 1;dino_sprite[2][94][7] = 1;dino_sprite[2][94][8] = 1;dino_sprite[2][94][9] = 1;dino_sprite[2][94][10] = 1;dino_sprite[2][94][11] = 1;dino_sprite[2][94][12] = 1;dino_sprite[2][94][13] = 1;dino_sprite[2][94][14] = 1;dino_sprite[2][94][15] = 1;dino_sprite[2][94][16] = 1;dino_sprite[2][94][17] = 1;dino_sprite[2][94][18] = 1;dino_sprite[2][94][19] = 1;dino_sprite[2][94][20] = 1;dino_sprite[2][94][21] = 1;dino_sprite[2][94][22] = 1;dino_sprite[2][94][23] = 1;dino_sprite[2][94][24] = 1;dino_sprite[2][94][25] = 1;dino_sprite[2][95][0] = 1;dino_sprite[2][95][1] = 1;dino_sprite[2][95][2] = 1;dino_sprite[2][95][3] = 1;dino_sprite[2][95][4] = 1;dino_sprite[2][95][5] = 1;dino_sprite[2][95][6] = 1;dino_sprite[2][95][7] = 1;dino_sprite[2][95][8] = 1;dino_sprite[2][95][9] = 1;dino_sprite[2][95][10] = 1;dino_sprite[2][95][11] = 1;dino_sprite[2][95][12] = 1;dino_sprite[2][95][13] = 1;dino_sprite[2][95][14] = 1;dino_sprite[2][95][15] = 1;dino_sprite[2][95][16] = 1;dino_sprite[2][95][17] = 1;dino_sprite[2][95][18] = 1;dino_sprite[2][95][19] = 1;dino_sprite[2][95][20] = 1;dino_sprite[2][95][21] = 1;dino_sprite[2][95][22] = 1;dino_sprite[2][95][23] = 1;dino_sprite[2][95][24] = 1;dino_sprite[2][95][25] = 1;dino_sprite[2][96][3] = 1;dino_sprite[2][96][4] = 1;dino_sprite[2][96][5] = 1;dino_sprite[2][96][6] = 1;dino_sprite[2][96][7] = 1;dino_sprite[2][96][8] = 1;dino_sprite[2][96][9] = 1;dino_sprite[2][96][10] = 1;dino_sprite[2][96][11] = 1;dino_sprite[2][96][12] = 1;dino_sprite[2][96][13] = 1;dino_sprite[2][96][14] = 1;dino_sprite[2][96][15] = 1;dino_sprite[2][96][16] = 1;dino_sprite[2][96][17] = 1;dino_sprite[2][96][18] = 1;dino_sprite[2][96][19] = 1;dino_sprite[2][96][20] = 1;dino_sprite[2][96][21] = 1;dino_sprite[2][96][22] = 1;dino_sprite[2][96][23] = 1;dino_sprite[2][96][24] = 1;dino_sprite[2][96][25] = 1;dino_sprite[2][97][3] = 1;dino_sprite[2][97][4] = 1;dino_sprite[2][97][5] = 1;dino_sprite[2][97][6] = 1;dino_sprite[2][97][7] = 1;dino_sprite[2][97][8] = 1;dino_sprite[2][97][9] = 1;dino_sprite[2][97][10] = 1;dino_sprite[2][97][11] = 1;dino_sprite[2][97][12] = 1;dino_sprite[2][97][13] = 1;dino_sprite[2][97][14] = 1;dino_sprite[2][97][15] = 1;dino_sprite[2][97][16] = 1;dino_sprite[2][97][17] = 1;dino_sprite[2][97][18] = 1;dino_sprite[2][97][19] = 1;dino_sprite[2][97][20] = 1;dino_sprite[2][97][21] = 1;dino_sprite[2][97][22] = 1;dino_sprite[2][97][23] = 1;dino_sprite[2][97][24] = 1;dino_sprite[2][97][25] = 1;dino_sprite[2][98][3] = 1;dino_sprite[2][98][4] = 1;dino_sprite[2][98][5] = 1;dino_sprite[2][98][6] = 1;dino_sprite[2][98][7] = 1;dino_sprite[2][98][8] = 1;dino_sprite[2][98][9] = 1;dino_sprite[2][98][10] = 1;dino_sprite[2][98][11] = 1;dino_sprite[2][98][12] = 1;dino_sprite[2][98][13] = 1;dino_sprite[2][98][14] = 1;dino_sprite[2][98][15] = 1;dino_sprite[2][98][16] = 1;dino_sprite[2][98][17] = 1;dino_sprite[2][98][18] = 1;dino_sprite[2][98][19] = 1;dino_sprite[2][98][20] = 1;dino_sprite[2][98][21] = 1;dino_sprite[2][98][22] = 1;dino_sprite[2][98][23] = 1;dino_sprite[2][98][24] = 1;dino_sprite[2][98][25] = 1;
  
	
	if (dino_count == 5000000)
	begin
		dino_count = 0;
		if (dino_sprite_choice == 1)
			dino_sprite_choice = 2;
		else
			dino_sprite_choice = 1;
	end
		
	dino_count = dino_count + 1; 
	
	if (jump_chn > 0)
		dino_sprite_choice = 0; // JUMP
	
	
	if ((dyno_x >= 0 && dyno_x < 100) && (dyno_y >= 0 && dyno_y < 100)) begin
		if (dino_sprite[dino_sprite_choice][dyno_x][dyno_y] == 1) begin
			r = 1;
			g = 1;
			b = 1;
		end
	end
	
	
	// -- CACTUS_SPRITE_CHOICE --
	cactuses_sprite_choice[0] = 0; cactuses_sprite_choice[1] = 3; cactuses_sprite_choice[2] = 1; cactuses_sprite_choice[3] = 2; cactuses_sprite_choice[4] = 4; cactuses_sprite_choice[5] = 0; cactuses_sprite_choice[6] = 4; cactuses_sprite_choice[7] = 2; cactuses_sprite_choice[8] = 6; cactuses_sprite_choice[9] = 0; cactuses_sprite_choice[10] = 3; cactuses_sprite_choice[11] = 5; cactuses_sprite_choice[12] = 2; cactuses_sprite_choice[13] = 1; cactuses_sprite_choice[14] = 6; cactuses_sprite_choice[15] = 4; cactuses_sprite_choice[16] = 2; cactuses_sprite_choice[17] = 0; cactuses_sprite_choice[18] = 4; cactuses_sprite_choice[19] = 5; cactuses_sprite_choice[20] = 6; cactuses_sprite_choice[21] = 1; cactuses_sprite_choice[22] = 2; cactuses_sprite_choice[23] = 5; cactuses_sprite_choice[24] = 0; cactuses_sprite_choice[25] = 6; cactuses_sprite_choice[26] = 3; cactuses_sprite_choice[27] = 0; cactuses_sprite_choice[28] = 1; cactuses_sprite_choice[29] = 0; cactuses_sprite_choice[30] = 2; cactuses_sprite_choice[31] = 5;
	// -- CACTUS SPRITE --
	cactus_sprite[0][2][20] = 1;cactus_sprite[0][2][21] = 1;cactus_sprite[0][2][22] = 1;cactus_sprite[0][2][23] = 1;cactus_sprite[0][2][24] = 1;cactus_sprite[0][2][25] = 1;cactus_sprite[0][2][26] = 1;cactus_sprite[0][2][27] = 1;cactus_sprite[0][2][28] = 1;cactus_sprite[0][2][29] = 1;cactus_sprite[0][2][30] = 1;cactus_sprite[0][2][31] = 1;cactus_sprite[0][2][32] = 1;cactus_sprite[0][2][33] = 1;cactus_sprite[0][2][34] = 1;cactus_sprite[0][2][35] = 1;cactus_sprite[0][2][36] = 1;cactus_sprite[0][2][37] = 1;cactus_sprite[0][2][38] = 1;cactus_sprite[0][2][39] = 1;cactus_sprite[0][2][40] = 1;cactus_sprite[0][2][41] = 1;cactus_sprite[0][2][42] = 1;cactus_sprite[0][2][43] = 1;cactus_sprite[0][2][44] = 1;cactus_sprite[0][2][45] = 1;cactus_sprite[0][2][46] = 1;cactus_sprite[0][2][47] = 1;cactus_sprite[0][2][48] = 1;cactus_sprite[0][2][49] = 1;cactus_sprite[0][3][20] = 1;cactus_sprite[0][3][21] = 1;cactus_sprite[0][3][22] = 1;cactus_sprite[0][3][23] = 1;cactus_sprite[0][3][24] = 1;cactus_sprite[0][3][25] = 1;cactus_sprite[0][3][26] = 1;cactus_sprite[0][3][27] = 1;cactus_sprite[0][3][28] = 1;cactus_sprite[0][3][29] = 1;cactus_sprite[0][3][30] = 1;cactus_sprite[0][3][31] = 1;cactus_sprite[0][3][32] = 1;cactus_sprite[0][3][33] = 1;cactus_sprite[0][3][34] = 1;cactus_sprite[0][3][35] = 1;cactus_sprite[0][3][36] = 1;cactus_sprite[0][3][37] = 1;cactus_sprite[0][3][38] = 1;cactus_sprite[0][3][39] = 1;cactus_sprite[0][3][40] = 1;cactus_sprite[0][3][41] = 1;cactus_sprite[0][3][42] = 1;cactus_sprite[0][3][43] = 1;cactus_sprite[0][3][44] = 1;cactus_sprite[0][3][45] = 1;cactus_sprite[0][3][46] = 1;cactus_sprite[0][3][47] = 1;cactus_sprite[0][3][48] = 1;cactus_sprite[0][3][49] = 1;cactus_sprite[0][4][18] = 1;cactus_sprite[0][4][19] = 1;cactus_sprite[0][4][20] = 1;cactus_sprite[0][4][21] = 1;cactus_sprite[0][4][22] = 1;cactus_sprite[0][4][23] = 1;cactus_sprite[0][4][24] = 1;cactus_sprite[0][4][25] = 1;cactus_sprite[0][4][26] = 1;cactus_sprite[0][4][27] = 1;cactus_sprite[0][4][28] = 1;cactus_sprite[0][4][29] = 1;cactus_sprite[0][4][30] = 1;cactus_sprite[0][4][31] = 1;cactus_sprite[0][4][32] = 1;cactus_sprite[0][4][33] = 1;cactus_sprite[0][4][34] = 1;cactus_sprite[0][4][35] = 1;cactus_sprite[0][4][36] = 1;cactus_sprite[0][4][37] = 1;cactus_sprite[0][4][38] = 1;cactus_sprite[0][4][39] = 1;cactus_sprite[0][4][40] = 1;cactus_sprite[0][4][41] = 1;cactus_sprite[0][4][42] = 1;cactus_sprite[0][4][43] = 1;cactus_sprite[0][4][44] = 1;cactus_sprite[0][4][45] = 1;cactus_sprite[0][4][46] = 1;cactus_sprite[0][4][47] = 1;cactus_sprite[0][4][48] = 1;cactus_sprite[0][4][49] = 1;cactus_sprite[0][4][50] = 1;cactus_sprite[0][4][51] = 1;cactus_sprite[0][5][18] = 1;cactus_sprite[0][5][19] = 1;cactus_sprite[0][5][20] = 1;cactus_sprite[0][5][21] = 1;cactus_sprite[0][5][22] = 1;cactus_sprite[0][5][23] = 1;cactus_sprite[0][5][24] = 1;cactus_sprite[0][5][25] = 1;cactus_sprite[0][5][26] = 1;cactus_sprite[0][5][27] = 1;cactus_sprite[0][5][28] = 1;cactus_sprite[0][5][29] = 1;cactus_sprite[0][5][30] = 1;cactus_sprite[0][5][31] = 1;cactus_sprite[0][5][32] = 1;cactus_sprite[0][5][33] = 1;cactus_sprite[0][5][34] = 1;cactus_sprite[0][5][35] = 1;cactus_sprite[0][5][36] = 1;cactus_sprite[0][5][37] = 1;cactus_sprite[0][5][38] = 1;cactus_sprite[0][5][39] = 1;cactus_sprite[0][5][40] = 1;cactus_sprite[0][5][41] = 1;cactus_sprite[0][5][42] = 1;cactus_sprite[0][5][43] = 1;cactus_sprite[0][5][44] = 1;cactus_sprite[0][5][45] = 1;cactus_sprite[0][5][46] = 1;cactus_sprite[0][5][47] = 1;cactus_sprite[0][5][48] = 1;cactus_sprite[0][5][49] = 1;cactus_sprite[0][5][50] = 1;cactus_sprite[0][5][51] = 1;cactus_sprite[0][6][18] = 1;cactus_sprite[0][6][19] = 1;cactus_sprite[0][6][20] = 1;cactus_sprite[0][6][21] = 1;cactus_sprite[0][6][22] = 1;cactus_sprite[0][6][23] = 1;cactus_sprite[0][6][24] = 1;cactus_sprite[0][6][25] = 1;cactus_sprite[0][6][26] = 1;cactus_sprite[0][6][27] = 1;cactus_sprite[0][6][28] = 1;cactus_sprite[0][6][29] = 1;cactus_sprite[0][6][30] = 1;cactus_sprite[0][6][31] = 1;cactus_sprite[0][6][32] = 1;cactus_sprite[0][6][33] = 1;cactus_sprite[0][6][34] = 1;cactus_sprite[0][6][35] = 1;cactus_sprite[0][6][36] = 1;cactus_sprite[0][6][37] = 1;cactus_sprite[0][6][38] = 1;cactus_sprite[0][6][39] = 1;cactus_sprite[0][6][40] = 1;cactus_sprite[0][6][41] = 1;cactus_sprite[0][6][42] = 1;cactus_sprite[0][6][43] = 1;cactus_sprite[0][6][44] = 1;cactus_sprite[0][6][45] = 1;cactus_sprite[0][6][46] = 1;cactus_sprite[0][6][47] = 1;cactus_sprite[0][6][48] = 1;cactus_sprite[0][6][49] = 1;cactus_sprite[0][6][50] = 1;cactus_sprite[0][6][51] = 1;cactus_sprite[0][6][52] = 1;cactus_sprite[0][6][53] = 1;cactus_sprite[0][7][18] = 1;cactus_sprite[0][7][19] = 1;cactus_sprite[0][7][20] = 1;cactus_sprite[0][7][21] = 1;cactus_sprite[0][7][22] = 1;cactus_sprite[0][7][23] = 1;cactus_sprite[0][7][24] = 1;cactus_sprite[0][7][25] = 1;cactus_sprite[0][7][26] = 1;cactus_sprite[0][7][27] = 1;cactus_sprite[0][7][28] = 1;cactus_sprite[0][7][29] = 1;cactus_sprite[0][7][30] = 1;cactus_sprite[0][7][31] = 1;cactus_sprite[0][7][32] = 1;cactus_sprite[0][7][33] = 1;cactus_sprite[0][7][34] = 1;cactus_sprite[0][7][35] = 1;cactus_sprite[0][7][36] = 1;cactus_sprite[0][7][37] = 1;cactus_sprite[0][7][38] = 1;cactus_sprite[0][7][39] = 1;cactus_sprite[0][7][40] = 1;cactus_sprite[0][7][41] = 1;cactus_sprite[0][7][42] = 1;cactus_sprite[0][7][43] = 1;cactus_sprite[0][7][44] = 1;cactus_sprite[0][7][45] = 1;cactus_sprite[0][7][46] = 1;cactus_sprite[0][7][47] = 1;cactus_sprite[0][7][48] = 1;cactus_sprite[0][7][49] = 1;cactus_sprite[0][7][50] = 1;cactus_sprite[0][7][51] = 1;cactus_sprite[0][7][52] = 1;cactus_sprite[0][7][53] = 1;cactus_sprite[0][8][18] = 1;cactus_sprite[0][8][19] = 1;cactus_sprite[0][8][20] = 1;cactus_sprite[0][8][21] = 1;cactus_sprite[0][8][22] = 1;cactus_sprite[0][8][23] = 1;cactus_sprite[0][8][24] = 1;cactus_sprite[0][8][25] = 1;cactus_sprite[0][8][26] = 1;cactus_sprite[0][8][27] = 1;cactus_sprite[0][8][28] = 1;cactus_sprite[0][8][29] = 1;cactus_sprite[0][8][30] = 1;cactus_sprite[0][8][31] = 1;cactus_sprite[0][8][32] = 1;cactus_sprite[0][8][33] = 1;cactus_sprite[0][8][34] = 1;cactus_sprite[0][8][35] = 1;cactus_sprite[0][8][36] = 1;cactus_sprite[0][8][37] = 1;cactus_sprite[0][8][38] = 1;cactus_sprite[0][8][39] = 1;cactus_sprite[0][8][40] = 1;cactus_sprite[0][8][41] = 1;cactus_sprite[0][8][42] = 1;cactus_sprite[0][8][43] = 1;cactus_sprite[0][8][44] = 1;cactus_sprite[0][8][45] = 1;cactus_sprite[0][8][46] = 1;cactus_sprite[0][8][47] = 1;cactus_sprite[0][8][48] = 1;cactus_sprite[0][8][49] = 1;cactus_sprite[0][8][50] = 1;cactus_sprite[0][8][51] = 1;cactus_sprite[0][8][52] = 1;cactus_sprite[0][8][53] = 1;cactus_sprite[0][8][54] = 1;cactus_sprite[0][8][55] = 1;cactus_sprite[0][9][18] = 1;cactus_sprite[0][9][19] = 1;cactus_sprite[0][9][20] = 1;cactus_sprite[0][9][21] = 1;cactus_sprite[0][9][22] = 1;cactus_sprite[0][9][23] = 1;cactus_sprite[0][9][24] = 1;cactus_sprite[0][9][25] = 1;cactus_sprite[0][9][26] = 1;cactus_sprite[0][9][27] = 1;cactus_sprite[0][9][28] = 1;cactus_sprite[0][9][29] = 1;cactus_sprite[0][9][30] = 1;cactus_sprite[0][9][31] = 1;cactus_sprite[0][9][32] = 1;cactus_sprite[0][9][33] = 1;cactus_sprite[0][9][34] = 1;cactus_sprite[0][9][35] = 1;cactus_sprite[0][9][36] = 1;cactus_sprite[0][9][37] = 1;cactus_sprite[0][9][38] = 1;cactus_sprite[0][9][39] = 1;cactus_sprite[0][9][40] = 1;cactus_sprite[0][9][41] = 1;cactus_sprite[0][9][42] = 1;cactus_sprite[0][9][43] = 1;cactus_sprite[0][9][44] = 1;cactus_sprite[0][9][45] = 1;cactus_sprite[0][9][46] = 1;cactus_sprite[0][9][47] = 1;cactus_sprite[0][9][48] = 1;cactus_sprite[0][9][49] = 1;cactus_sprite[0][9][50] = 1;cactus_sprite[0][9][51] = 1;cactus_sprite[0][9][52] = 1;cactus_sprite[0][9][53] = 1;cactus_sprite[0][9][54] = 1;cactus_sprite[0][9][55] = 1;cactus_sprite[0][10][20] = 1;cactus_sprite[0][10][21] = 1;cactus_sprite[0][10][22] = 1;cactus_sprite[0][10][23] = 1;cactus_sprite[0][10][24] = 1;cactus_sprite[0][10][25] = 1;cactus_sprite[0][10][26] = 1;cactus_sprite[0][10][27] = 1;cactus_sprite[0][10][28] = 1;cactus_sprite[0][10][29] = 1;cactus_sprite[0][10][30] = 1;cactus_sprite[0][10][31] = 1;cactus_sprite[0][10][32] = 1;cactus_sprite[0][10][33] = 1;cactus_sprite[0][10][34] = 1;cactus_sprite[0][10][35] = 1;cactus_sprite[0][10][36] = 1;cactus_sprite[0][10][37] = 1;cactus_sprite[0][10][38] = 1;cactus_sprite[0][10][39] = 1;cactus_sprite[0][10][40] = 1;cactus_sprite[0][10][41] = 1;cactus_sprite[0][10][42] = 1;cactus_sprite[0][10][43] = 1;cactus_sprite[0][10][44] = 1;cactus_sprite[0][10][45] = 1;cactus_sprite[0][10][46] = 1;cactus_sprite[0][10][47] = 1;cactus_sprite[0][10][48] = 1;cactus_sprite[0][10][49] = 1;cactus_sprite[0][10][50] = 1;cactus_sprite[0][10][51] = 1;cactus_sprite[0][10][52] = 1;cactus_sprite[0][10][53] = 1;cactus_sprite[0][10][54] = 1;cactus_sprite[0][10][55] = 1;cactus_sprite[0][10][56] = 1;cactus_sprite[0][10][57] = 1;cactus_sprite[0][11][20] = 1;cactus_sprite[0][11][21] = 1;cactus_sprite[0][11][22] = 1;cactus_sprite[0][11][23] = 1;cactus_sprite[0][11][24] = 1;cactus_sprite[0][11][25] = 1;cactus_sprite[0][11][26] = 1;cactus_sprite[0][11][27] = 1;cactus_sprite[0][11][28] = 1;cactus_sprite[0][11][29] = 1;cactus_sprite[0][11][30] = 1;cactus_sprite[0][11][31] = 1;cactus_sprite[0][11][32] = 1;cactus_sprite[0][11][33] = 1;cactus_sprite[0][11][34] = 1;cactus_sprite[0][11][35] = 1;cactus_sprite[0][11][36] = 1;cactus_sprite[0][11][37] = 1;cactus_sprite[0][11][38] = 1;cactus_sprite[0][11][39] = 1;cactus_sprite[0][11][40] = 1;cactus_sprite[0][11][41] = 1;cactus_sprite[0][11][42] = 1;cactus_sprite[0][11][43] = 1;cactus_sprite[0][11][44] = 1;cactus_sprite[0][11][45] = 1;cactus_sprite[0][11][46] = 1;cactus_sprite[0][11][47] = 1;cactus_sprite[0][11][48] = 1;cactus_sprite[0][11][49] = 1;cactus_sprite[0][11][50] = 1;cactus_sprite[0][11][51] = 1;cactus_sprite[0][11][52] = 1;cactus_sprite[0][11][53] = 1;cactus_sprite[0][11][54] = 1;cactus_sprite[0][11][55] = 1;cactus_sprite[0][11][56] = 1;cactus_sprite[0][11][57] = 1;cactus_sprite[0][12][48] = 1;cactus_sprite[0][12][49] = 1;cactus_sprite[0][12][50] = 1;cactus_sprite[0][12][51] = 1;cactus_sprite[0][12][52] = 1;cactus_sprite[0][12][53] = 1;cactus_sprite[0][12][54] = 1;cactus_sprite[0][12][55] = 1;cactus_sprite[0][12][56] = 1;cactus_sprite[0][12][57] = 1;cactus_sprite[0][13][48] = 1;cactus_sprite[0][13][49] = 1;cactus_sprite[0][13][50] = 1;cactus_sprite[0][13][51] = 1;cactus_sprite[0][13][52] = 1;cactus_sprite[0][13][53] = 1;cactus_sprite[0][13][54] = 1;cactus_sprite[0][13][55] = 1;cactus_sprite[0][13][56] = 1;cactus_sprite[0][13][57] = 1;cactus_sprite[0][14][48] = 1;cactus_sprite[0][14][49] = 1;cactus_sprite[0][14][50] = 1;cactus_sprite[0][14][51] = 1;cactus_sprite[0][14][52] = 1;cactus_sprite[0][14][53] = 1;cactus_sprite[0][14][54] = 1;cactus_sprite[0][14][55] = 1;cactus_sprite[0][14][56] = 1;cactus_sprite[0][14][57] = 1;cactus_sprite[0][15][48] = 1;cactus_sprite[0][15][49] = 1;cactus_sprite[0][15][50] = 1;cactus_sprite[0][15][51] = 1;cactus_sprite[0][15][52] = 1;cactus_sprite[0][15][53] = 1;cactus_sprite[0][15][54] = 1;cactus_sprite[0][15][55] = 1;cactus_sprite[0][15][56] = 1;cactus_sprite[0][15][57] = 1;cactus_sprite[0][16][48] = 1;cactus_sprite[0][16][49] = 1;cactus_sprite[0][16][50] = 1;cactus_sprite[0][16][51] = 1;cactus_sprite[0][16][52] = 1;cactus_sprite[0][16][53] = 1;cactus_sprite[0][16][54] = 1;cactus_sprite[0][16][55] = 1;cactus_sprite[0][16][56] = 1;cactus_sprite[0][16][57] = 1;cactus_sprite[0][17][48] = 1;cactus_sprite[0][17][49] = 1;cactus_sprite[0][17][50] = 1;cactus_sprite[0][17][51] = 1;cactus_sprite[0][17][52] = 1;cactus_sprite[0][17][53] = 1;cactus_sprite[0][17][54] = 1;cactus_sprite[0][17][55] = 1;cactus_sprite[0][17][56] = 1;cactus_sprite[0][17][57] = 1;cactus_sprite[0][18][10] = 1;cactus_sprite[0][18][11] = 1;cactus_sprite[0][18][12] = 1;cactus_sprite[0][18][13] = 1;cactus_sprite[0][18][14] = 1;cactus_sprite[0][18][15] = 1;cactus_sprite[0][18][16] = 1;cactus_sprite[0][18][17] = 1;cactus_sprite[0][18][18] = 1;cactus_sprite[0][18][19] = 1;cactus_sprite[0][18][20] = 1;cactus_sprite[0][18][21] = 1;cactus_sprite[0][18][22] = 1;cactus_sprite[0][18][23] = 1;cactus_sprite[0][18][24] = 1;cactus_sprite[0][18][25] = 1;cactus_sprite[0][18][26] = 1;cactus_sprite[0][18][27] = 1;cactus_sprite[0][18][28] = 1;cactus_sprite[0][18][29] = 1;cactus_sprite[0][18][30] = 1;cactus_sprite[0][18][31] = 1;cactus_sprite[0][18][32] = 1;cactus_sprite[0][18][33] = 1;cactus_sprite[0][18][34] = 1;cactus_sprite[0][18][35] = 1;cactus_sprite[0][18][36] = 1;cactus_sprite[0][18][37] = 1;cactus_sprite[0][18][38] = 1;cactus_sprite[0][18][39] = 1;cactus_sprite[0][18][40] = 1;cactus_sprite[0][18][41] = 1;cactus_sprite[0][18][42] = 1;cactus_sprite[0][18][43] = 1;cactus_sprite[0][18][44] = 1;cactus_sprite[0][18][45] = 1;cactus_sprite[0][18][46] = 1;cactus_sprite[0][18][47] = 1;cactus_sprite[0][18][48] = 1;cactus_sprite[0][18][49] = 1;cactus_sprite[0][18][50] = 1;cactus_sprite[0][18][51] = 1;cactus_sprite[0][18][52] = 1;cactus_sprite[0][18][53] = 1;cactus_sprite[0][18][54] = 1;cactus_sprite[0][18][55] = 1;cactus_sprite[0][18][56] = 1;cactus_sprite[0][18][57] = 1;cactus_sprite[0][18][58] = 1;cactus_sprite[0][18][59] = 1;cactus_sprite[0][18][60] = 1;cactus_sprite[0][18][61] = 1;cactus_sprite[0][18][62] = 1;cactus_sprite[0][18][63] = 1;cactus_sprite[0][18][64] = 1;cactus_sprite[0][18][65] = 1;cactus_sprite[0][18][66] = 1;cactus_sprite[0][18][67] = 1;cactus_sprite[0][18][68] = 1;cactus_sprite[0][18][69] = 1;cactus_sprite[0][18][70] = 1;cactus_sprite[0][18][71] = 1;cactus_sprite[0][18][72] = 1;cactus_sprite[0][18][73] = 1;cactus_sprite[0][18][74] = 1;cactus_sprite[0][18][75] = 1;cactus_sprite[0][18][76] = 1;cactus_sprite[0][18][77] = 1;cactus_sprite[0][18][78] = 1;cactus_sprite[0][18][79] = 1;cactus_sprite[0][18][80] = 1;cactus_sprite[0][18][81] = 1;cactus_sprite[0][18][82] = 1;cactus_sprite[0][18][83] = 1;cactus_sprite[0][18][84] = 1;cactus_sprite[0][18][85] = 1;cactus_sprite[0][18][86] = 1;cactus_sprite[0][18][87] = 1;cactus_sprite[0][18][88] = 1;cactus_sprite[0][18][89] = 1;cactus_sprite[0][18][90] = 1;cactus_sprite[0][18][91] = 1;cactus_sprite[0][18][92] = 1;cactus_sprite[0][18][93] = 1;cactus_sprite[0][18][94] = 1;cactus_sprite[0][18][95] = 1;cactus_sprite[0][18][96] = 1;cactus_sprite[0][18][97] = 1;cactus_sprite[0][18][98] = 1;cactus_sprite[0][18][99] = 1;cactus_sprite[0][19][10] = 1;cactus_sprite[0][19][11] = 1;cactus_sprite[0][19][12] = 1;cactus_sprite[0][19][13] = 1;cactus_sprite[0][19][14] = 1;cactus_sprite[0][19][15] = 1;cactus_sprite[0][19][16] = 1;cactus_sprite[0][19][17] = 1;cactus_sprite[0][19][18] = 1;cactus_sprite[0][19][19] = 1;cactus_sprite[0][19][20] = 1;cactus_sprite[0][19][21] = 1;cactus_sprite[0][19][22] = 1;cactus_sprite[0][19][23] = 1;cactus_sprite[0][19][24] = 1;cactus_sprite[0][19][25] = 1;cactus_sprite[0][19][26] = 1;cactus_sprite[0][19][27] = 1;cactus_sprite[0][19][28] = 1;cactus_sprite[0][19][29] = 1;cactus_sprite[0][19][30] = 1;cactus_sprite[0][19][31] = 1;cactus_sprite[0][19][32] = 1;cactus_sprite[0][19][33] = 1;cactus_sprite[0][19][34] = 1;cactus_sprite[0][19][35] = 1;cactus_sprite[0][19][36] = 1;cactus_sprite[0][19][37] = 1;cactus_sprite[0][19][38] = 1;cactus_sprite[0][19][39] = 1;cactus_sprite[0][19][40] = 1;cactus_sprite[0][19][41] = 1;cactus_sprite[0][19][42] = 1;cactus_sprite[0][19][43] = 1;cactus_sprite[0][19][44] = 1;cactus_sprite[0][19][45] = 1;cactus_sprite[0][19][46] = 1;cactus_sprite[0][19][47] = 1;cactus_sprite[0][19][48] = 1;cactus_sprite[0][19][49] = 1;cactus_sprite[0][19][50] = 1;cactus_sprite[0][19][51] = 1;cactus_sprite[0][19][52] = 1;cactus_sprite[0][19][53] = 1;cactus_sprite[0][19][54] = 1;cactus_sprite[0][19][55] = 1;cactus_sprite[0][19][56] = 1;cactus_sprite[0][19][57] = 1;cactus_sprite[0][19][58] = 1;cactus_sprite[0][19][59] = 1;cactus_sprite[0][19][60] = 1;cactus_sprite[0][19][61] = 1;cactus_sprite[0][19][62] = 1;cactus_sprite[0][19][63] = 1;cactus_sprite[0][19][64] = 1;cactus_sprite[0][19][65] = 1;cactus_sprite[0][19][66] = 1;cactus_sprite[0][19][67] = 1;cactus_sprite[0][19][68] = 1;cactus_sprite[0][19][69] = 1;cactus_sprite[0][19][70] = 1;cactus_sprite[0][19][71] = 1;cactus_sprite[0][19][72] = 1;cactus_sprite[0][19][73] = 1;cactus_sprite[0][19][74] = 1;cactus_sprite[0][19][75] = 1;cactus_sprite[0][19][76] = 1;cactus_sprite[0][19][77] = 1;cactus_sprite[0][19][78] = 1;cactus_sprite[0][19][79] = 1;cactus_sprite[0][19][80] = 1;cactus_sprite[0][19][81] = 1;cactus_sprite[0][19][82] = 1;cactus_sprite[0][19][83] = 1;cactus_sprite[0][19][84] = 1;cactus_sprite[0][19][85] = 1;cactus_sprite[0][19][86] = 1;cactus_sprite[0][19][87] = 1;cactus_sprite[0][19][88] = 1;cactus_sprite[0][19][89] = 1;cactus_sprite[0][19][90] = 1;cactus_sprite[0][19][91] = 1;cactus_sprite[0][19][92] = 1;cactus_sprite[0][19][93] = 1;cactus_sprite[0][19][94] = 1;cactus_sprite[0][19][95] = 1;cactus_sprite[0][19][96] = 1;cactus_sprite[0][19][97] = 1;cactus_sprite[0][19][98] = 1;cactus_sprite[0][19][99] = 1;cactus_sprite[0][20][8] = 1;cactus_sprite[0][20][9] = 1;cactus_sprite[0][20][10] = 1;cactus_sprite[0][20][11] = 1;cactus_sprite[0][20][12] = 1;cactus_sprite[0][20][13] = 1;cactus_sprite[0][20][14] = 1;cactus_sprite[0][20][15] = 1;cactus_sprite[0][20][16] = 1;cactus_sprite[0][20][17] = 1;cactus_sprite[0][20][18] = 1;cactus_sprite[0][20][19] = 1;cactus_sprite[0][20][20] = 1;cactus_sprite[0][20][21] = 1;cactus_sprite[0][20][22] = 1;cactus_sprite[0][20][23] = 1;cactus_sprite[0][20][24] = 1;cactus_sprite[0][20][25] = 1;cactus_sprite[0][20][26] = 1;cactus_sprite[0][20][27] = 1;cactus_sprite[0][20][28] = 1;cactus_sprite[0][20][29] = 1;cactus_sprite[0][20][30] = 1;cactus_sprite[0][20][31] = 1;cactus_sprite[0][20][32] = 1;cactus_sprite[0][20][33] = 1;cactus_sprite[0][20][34] = 1;cactus_sprite[0][20][35] = 1;cactus_sprite[0][20][36] = 1;cactus_sprite[0][20][37] = 1;cactus_sprite[0][20][38] = 1;cactus_sprite[0][20][39] = 1;cactus_sprite[0][20][40] = 1;cactus_sprite[0][20][41] = 1;cactus_sprite[0][20][42] = 1;cactus_sprite[0][20][43] = 1;cactus_sprite[0][20][44] = 1;cactus_sprite[0][20][45] = 1;cactus_sprite[0][20][46] = 1;cactus_sprite[0][20][47] = 1;cactus_sprite[0][20][48] = 1;cactus_sprite[0][20][49] = 1;cactus_sprite[0][20][50] = 1;cactus_sprite[0][20][51] = 1;cactus_sprite[0][20][52] = 1;cactus_sprite[0][20][53] = 1;cactus_sprite[0][20][54] = 1;cactus_sprite[0][20][55] = 1;cactus_sprite[0][20][56] = 1;cactus_sprite[0][20][57] = 1;cactus_sprite[0][20][58] = 1;cactus_sprite[0][20][59] = 1;cactus_sprite[0][20][60] = 1;cactus_sprite[0][20][61] = 1;cactus_sprite[0][20][62] = 1;cactus_sprite[0][20][63] = 1;cactus_sprite[0][20][64] = 1;cactus_sprite[0][20][65] = 1;cactus_sprite[0][20][66] = 1;cactus_sprite[0][20][67] = 1;cactus_sprite[0][20][68] = 1;cactus_sprite[0][20][69] = 1;cactus_sprite[0][20][70] = 1;cactus_sprite[0][20][71] = 1;cactus_sprite[0][20][72] = 1;cactus_sprite[0][20][73] = 1;cactus_sprite[0][20][74] = 1;cactus_sprite[0][20][75] = 1;cactus_sprite[0][20][76] = 1;cactus_sprite[0][20][77] = 1;cactus_sprite[0][20][78] = 1;cactus_sprite[0][20][79] = 1;cactus_sprite[0][20][80] = 1;cactus_sprite[0][20][81] = 1;cactus_sprite[0][20][82] = 1;cactus_sprite[0][20][83] = 1;cactus_sprite[0][20][84] = 1;cactus_sprite[0][20][85] = 1;cactus_sprite[0][20][86] = 1;cactus_sprite[0][20][87] = 1;cactus_sprite[0][20][88] = 1;cactus_sprite[0][20][89] = 1;cactus_sprite[0][20][90] = 1;cactus_sprite[0][20][91] = 1;cactus_sprite[0][20][92] = 1;cactus_sprite[0][20][93] = 1;cactus_sprite[0][20][94] = 1;cactus_sprite[0][20][95] = 1;cactus_sprite[0][20][96] = 1;cactus_sprite[0][20][97] = 1;cactus_sprite[0][20][98] = 1;cactus_sprite[0][20][99] = 1;cactus_sprite[0][21][8] = 1;cactus_sprite[0][21][9] = 1;cactus_sprite[0][21][10] = 1;cactus_sprite[0][21][11] = 1;cactus_sprite[0][21][12] = 1;cactus_sprite[0][21][13] = 1;cactus_sprite[0][21][14] = 1;cactus_sprite[0][21][15] = 1;cactus_sprite[0][21][16] = 1;cactus_sprite[0][21][17] = 1;cactus_sprite[0][21][18] = 1;cactus_sprite[0][21][19] = 1;cactus_sprite[0][21][20] = 1;cactus_sprite[0][21][21] = 1;cactus_sprite[0][21][22] = 1;cactus_sprite[0][21][23] = 1;cactus_sprite[0][21][24] = 1;cactus_sprite[0][21][25] = 1;cactus_sprite[0][21][26] = 1;cactus_sprite[0][21][27] = 1;cactus_sprite[0][21][28] = 1;cactus_sprite[0][21][29] = 1;cactus_sprite[0][21][30] = 1;cactus_sprite[0][21][31] = 1;cactus_sprite[0][21][32] = 1;cactus_sprite[0][21][33] = 1;cactus_sprite[0][21][34] = 1;cactus_sprite[0][21][35] = 1;cactus_sprite[0][21][36] = 1;cactus_sprite[0][21][37] = 1;cactus_sprite[0][21][38] = 1;cactus_sprite[0][21][39] = 1;cactus_sprite[0][21][40] = 1;cactus_sprite[0][21][41] = 1;cactus_sprite[0][21][42] = 1;cactus_sprite[0][21][43] = 1;cactus_sprite[0][21][44] = 1;cactus_sprite[0][21][45] = 1;cactus_sprite[0][21][46] = 1;cactus_sprite[0][21][47] = 1;cactus_sprite[0][21][48] = 1;cactus_sprite[0][21][49] = 1;cactus_sprite[0][21][50] = 1;cactus_sprite[0][21][51] = 1;cactus_sprite[0][21][52] = 1;cactus_sprite[0][21][53] = 1;cactus_sprite[0][21][54] = 1;cactus_sprite[0][21][55] = 1;cactus_sprite[0][21][56] = 1;cactus_sprite[0][21][57] = 1;cactus_sprite[0][21][58] = 1;cactus_sprite[0][21][59] = 1;cactus_sprite[0][21][60] = 1;cactus_sprite[0][21][61] = 1;cactus_sprite[0][21][62] = 1;cactus_sprite[0][21][63] = 1;cactus_sprite[0][21][64] = 1;cactus_sprite[0][21][65] = 1;cactus_sprite[0][21][66] = 1;cactus_sprite[0][21][67] = 1;cactus_sprite[0][21][68] = 1;cactus_sprite[0][21][69] = 1;cactus_sprite[0][21][70] = 1;cactus_sprite[0][21][71] = 1;cactus_sprite[0][21][72] = 1;cactus_sprite[0][21][73] = 1;cactus_sprite[0][21][74] = 1;cactus_sprite[0][21][75] = 1;cactus_sprite[0][21][76] = 1;cactus_sprite[0][21][77] = 1;cactus_sprite[0][21][78] = 1;cactus_sprite[0][21][79] = 1;cactus_sprite[0][21][80] = 1;cactus_sprite[0][21][81] = 1;cactus_sprite[0][21][82] = 1;cactus_sprite[0][21][83] = 1;cactus_sprite[0][21][84] = 1;cactus_sprite[0][21][85] = 1;cactus_sprite[0][21][86] = 1;cactus_sprite[0][21][87] = 1;cactus_sprite[0][21][88] = 1;cactus_sprite[0][21][89] = 1;cactus_sprite[0][21][90] = 1;cactus_sprite[0][21][91] = 1;cactus_sprite[0][21][92] = 1;cactus_sprite[0][21][93] = 1;cactus_sprite[0][21][94] = 1;cactus_sprite[0][21][95] = 1;cactus_sprite[0][21][96] = 1;cactus_sprite[0][21][97] = 1;cactus_sprite[0][21][98] = 1;cactus_sprite[0][21][99] = 1;cactus_sprite[0][22][8] = 1;cactus_sprite[0][22][9] = 1;cactus_sprite[0][22][10] = 1;cactus_sprite[0][22][11] = 1;cactus_sprite[0][22][12] = 1;cactus_sprite[0][22][13] = 1;cactus_sprite[0][22][14] = 1;cactus_sprite[0][22][15] = 1;cactus_sprite[0][22][16] = 1;cactus_sprite[0][22][17] = 1;cactus_sprite[0][22][18] = 1;cactus_sprite[0][22][19] = 1;cactus_sprite[0][22][20] = 1;cactus_sprite[0][22][21] = 1;cactus_sprite[0][22][22] = 1;cactus_sprite[0][22][23] = 1;cactus_sprite[0][22][24] = 1;cactus_sprite[0][22][25] = 1;cactus_sprite[0][22][26] = 1;cactus_sprite[0][22][27] = 1;cactus_sprite[0][22][28] = 1;cactus_sprite[0][22][29] = 1;cactus_sprite[0][22][30] = 1;cactus_sprite[0][22][31] = 1;cactus_sprite[0][22][32] = 1;cactus_sprite[0][22][33] = 1;cactus_sprite[0][22][34] = 1;cactus_sprite[0][22][35] = 1;cactus_sprite[0][22][36] = 1;cactus_sprite[0][22][37] = 1;cactus_sprite[0][22][38] = 1;cactus_sprite[0][22][39] = 1;cactus_sprite[0][22][40] = 1;cactus_sprite[0][22][41] = 1;cactus_sprite[0][22][42] = 1;cactus_sprite[0][22][43] = 1;cactus_sprite[0][22][44] = 1;cactus_sprite[0][22][45] = 1;cactus_sprite[0][22][46] = 1;cactus_sprite[0][22][47] = 1;cactus_sprite[0][22][48] = 1;cactus_sprite[0][22][49] = 1;cactus_sprite[0][22][50] = 1;cactus_sprite[0][22][51] = 1;cactus_sprite[0][22][52] = 1;cactus_sprite[0][22][53] = 1;cactus_sprite[0][22][54] = 1;cactus_sprite[0][22][55] = 1;cactus_sprite[0][22][56] = 1;cactus_sprite[0][22][57] = 1;cactus_sprite[0][22][58] = 1;cactus_sprite[0][22][59] = 1;cactus_sprite[0][22][60] = 1;cactus_sprite[0][22][61] = 1;cactus_sprite[0][22][62] = 1;cactus_sprite[0][22][63] = 1;cactus_sprite[0][22][64] = 1;cactus_sprite[0][22][65] = 1;cactus_sprite[0][22][66] = 1;cactus_sprite[0][22][67] = 1;cactus_sprite[0][22][68] = 1;cactus_sprite[0][22][69] = 1;cactus_sprite[0][22][70] = 1;cactus_sprite[0][22][71] = 1;cactus_sprite[0][22][72] = 1;cactus_sprite[0][22][73] = 1;cactus_sprite[0][22][74] = 1;cactus_sprite[0][22][75] = 1;cactus_sprite[0][22][76] = 1;cactus_sprite[0][22][77] = 1;cactus_sprite[0][22][78] = 1;cactus_sprite[0][22][79] = 1;cactus_sprite[0][22][80] = 1;cactus_sprite[0][22][81] = 1;cactus_sprite[0][22][82] = 1;cactus_sprite[0][22][83] = 1;cactus_sprite[0][22][84] = 1;cactus_sprite[0][22][85] = 1;cactus_sprite[0][22][86] = 1;cactus_sprite[0][22][87] = 1;cactus_sprite[0][22][88] = 1;cactus_sprite[0][22][89] = 1;cactus_sprite[0][22][90] = 1;cactus_sprite[0][22][91] = 1;cactus_sprite[0][22][92] = 1;cactus_sprite[0][22][93] = 1;cactus_sprite[0][22][94] = 1;cactus_sprite[0][22][95] = 1;cactus_sprite[0][22][96] = 1;cactus_sprite[0][22][97] = 1;cactus_sprite[0][22][98] = 1;cactus_sprite[0][22][99] = 1;cactus_sprite[0][23][8] = 1;cactus_sprite[0][23][9] = 1;cactus_sprite[0][23][10] = 1;cactus_sprite[0][23][11] = 1;cactus_sprite[0][23][12] = 1;cactus_sprite[0][23][13] = 1;cactus_sprite[0][23][14] = 1;cactus_sprite[0][23][15] = 1;cactus_sprite[0][23][16] = 1;cactus_sprite[0][23][17] = 1;cactus_sprite[0][23][18] = 1;cactus_sprite[0][23][19] = 1;cactus_sprite[0][23][20] = 1;cactus_sprite[0][23][21] = 1;cactus_sprite[0][23][22] = 1;cactus_sprite[0][23][23] = 1;cactus_sprite[0][23][24] = 1;cactus_sprite[0][23][25] = 1;cactus_sprite[0][23][26] = 1;cactus_sprite[0][23][27] = 1;cactus_sprite[0][23][28] = 1;cactus_sprite[0][23][29] = 1;cactus_sprite[0][23][30] = 1;cactus_sprite[0][23][31] = 1;cactus_sprite[0][23][32] = 1;cactus_sprite[0][23][33] = 1;cactus_sprite[0][23][34] = 1;cactus_sprite[0][23][35] = 1;cactus_sprite[0][23][36] = 1;cactus_sprite[0][23][37] = 1;cactus_sprite[0][23][38] = 1;cactus_sprite[0][23][39] = 1;cactus_sprite[0][23][40] = 1;cactus_sprite[0][23][41] = 1;cactus_sprite[0][23][42] = 1;cactus_sprite[0][23][43] = 1;cactus_sprite[0][23][44] = 1;cactus_sprite[0][23][45] = 1;cactus_sprite[0][23][46] = 1;cactus_sprite[0][23][47] = 1;cactus_sprite[0][23][48] = 1;cactus_sprite[0][23][49] = 1;cactus_sprite[0][23][50] = 1;cactus_sprite[0][23][51] = 1;cactus_sprite[0][23][52] = 1;cactus_sprite[0][23][53] = 1;cactus_sprite[0][23][54] = 1;cactus_sprite[0][23][55] = 1;cactus_sprite[0][23][56] = 1;cactus_sprite[0][23][57] = 1;cactus_sprite[0][23][58] = 1;cactus_sprite[0][23][59] = 1;cactus_sprite[0][23][60] = 1;cactus_sprite[0][23][61] = 1;cactus_sprite[0][23][62] = 1;cactus_sprite[0][23][63] = 1;cactus_sprite[0][23][64] = 1;cactus_sprite[0][23][65] = 1;cactus_sprite[0][23][66] = 1;cactus_sprite[0][23][67] = 1;cactus_sprite[0][23][68] = 1;cactus_sprite[0][23][69] = 1;cactus_sprite[0][23][70] = 1;cactus_sprite[0][23][71] = 1;cactus_sprite[0][23][72] = 1;cactus_sprite[0][23][73] = 1;cactus_sprite[0][23][74] = 1;cactus_sprite[0][23][75] = 1;cactus_sprite[0][23][76] = 1;cactus_sprite[0][23][77] = 1;cactus_sprite[0][23][78] = 1;cactus_sprite[0][23][79] = 1;cactus_sprite[0][23][80] = 1;cactus_sprite[0][23][81] = 1;cactus_sprite[0][23][82] = 1;cactus_sprite[0][23][83] = 1;cactus_sprite[0][23][84] = 1;cactus_sprite[0][23][85] = 1;cactus_sprite[0][23][86] = 1;cactus_sprite[0][23][87] = 1;cactus_sprite[0][23][88] = 1;cactus_sprite[0][23][89] = 1;cactus_sprite[0][23][90] = 1;cactus_sprite[0][23][91] = 1;cactus_sprite[0][23][92] = 1;cactus_sprite[0][23][93] = 1;cactus_sprite[0][23][94] = 1;cactus_sprite[0][23][95] = 1;cactus_sprite[0][23][96] = 1;cactus_sprite[0][23][97] = 1;cactus_sprite[0][23][98] = 1;cactus_sprite[0][23][99] = 1;cactus_sprite[0][24][8] = 1;cactus_sprite[0][24][9] = 1;cactus_sprite[0][24][10] = 1;cactus_sprite[0][24][11] = 1;cactus_sprite[0][24][12] = 1;cactus_sprite[0][24][13] = 1;cactus_sprite[0][24][14] = 1;cactus_sprite[0][24][15] = 1;cactus_sprite[0][24][16] = 1;cactus_sprite[0][24][17] = 1;cactus_sprite[0][24][18] = 1;cactus_sprite[0][24][19] = 1;cactus_sprite[0][24][20] = 1;cactus_sprite[0][24][21] = 1;cactus_sprite[0][24][22] = 1;cactus_sprite[0][24][23] = 1;cactus_sprite[0][24][24] = 1;cactus_sprite[0][24][25] = 1;cactus_sprite[0][24][26] = 1;cactus_sprite[0][24][27] = 1;cactus_sprite[0][24][28] = 1;cactus_sprite[0][24][29] = 1;cactus_sprite[0][24][30] = 1;cactus_sprite[0][24][31] = 1;cactus_sprite[0][24][32] = 1;cactus_sprite[0][24][33] = 1;cactus_sprite[0][24][34] = 1;cactus_sprite[0][24][35] = 1;cactus_sprite[0][24][36] = 1;cactus_sprite[0][24][37] = 1;cactus_sprite[0][24][38] = 1;cactus_sprite[0][24][39] = 1;cactus_sprite[0][24][40] = 1;cactus_sprite[0][24][41] = 1;cactus_sprite[0][24][42] = 1;cactus_sprite[0][24][43] = 1;cactus_sprite[0][24][44] = 1;cactus_sprite[0][24][45] = 1;cactus_sprite[0][24][46] = 1;cactus_sprite[0][24][47] = 1;cactus_sprite[0][24][48] = 1;cactus_sprite[0][24][49] = 1;cactus_sprite[0][24][50] = 1;cactus_sprite[0][24][51] = 1;cactus_sprite[0][24][52] = 1;cactus_sprite[0][24][53] = 1;cactus_sprite[0][24][54] = 1;cactus_sprite[0][24][55] = 1;cactus_sprite[0][24][56] = 1;cactus_sprite[0][24][57] = 1;cactus_sprite[0][24][58] = 1;cactus_sprite[0][24][59] = 1;cactus_sprite[0][24][60] = 1;cactus_sprite[0][24][61] = 1;cactus_sprite[0][24][62] = 1;cactus_sprite[0][24][63] = 1;cactus_sprite[0][24][64] = 1;cactus_sprite[0][24][65] = 1;cactus_sprite[0][24][66] = 1;cactus_sprite[0][24][67] = 1;cactus_sprite[0][24][68] = 1;cactus_sprite[0][24][69] = 1;cactus_sprite[0][24][70] = 1;cactus_sprite[0][24][71] = 1;cactus_sprite[0][24][72] = 1;cactus_sprite[0][24][73] = 1;cactus_sprite[0][24][74] = 1;cactus_sprite[0][24][75] = 1;cactus_sprite[0][24][76] = 1;cactus_sprite[0][24][77] = 1;cactus_sprite[0][24][78] = 1;cactus_sprite[0][24][79] = 1;cactus_sprite[0][24][80] = 1;cactus_sprite[0][24][81] = 1;cactus_sprite[0][24][82] = 1;cactus_sprite[0][24][83] = 1;cactus_sprite[0][24][84] = 1;cactus_sprite[0][24][85] = 1;cactus_sprite[0][24][86] = 1;cactus_sprite[0][24][87] = 1;cactus_sprite[0][24][88] = 1;cactus_sprite[0][24][89] = 1;cactus_sprite[0][24][90] = 1;cactus_sprite[0][24][91] = 1;cactus_sprite[0][24][92] = 1;cactus_sprite[0][24][93] = 1;cactus_sprite[0][24][94] = 1;cactus_sprite[0][24][95] = 1;cactus_sprite[0][24][96] = 1;cactus_sprite[0][24][97] = 1;cactus_sprite[0][24][98] = 1;cactus_sprite[0][24][99] = 1;cactus_sprite[0][25][8] = 1;cactus_sprite[0][25][9] = 1;cactus_sprite[0][25][10] = 1;cactus_sprite[0][25][11] = 1;cactus_sprite[0][25][12] = 1;cactus_sprite[0][25][13] = 1;cactus_sprite[0][25][14] = 1;cactus_sprite[0][25][15] = 1;cactus_sprite[0][25][16] = 1;cactus_sprite[0][25][17] = 1;cactus_sprite[0][25][18] = 1;cactus_sprite[0][25][19] = 1;cactus_sprite[0][25][20] = 1;cactus_sprite[0][25][21] = 1;cactus_sprite[0][25][22] = 1;cactus_sprite[0][25][23] = 1;cactus_sprite[0][25][24] = 1;cactus_sprite[0][25][25] = 1;cactus_sprite[0][25][26] = 1;cactus_sprite[0][25][27] = 1;cactus_sprite[0][25][28] = 1;cactus_sprite[0][25][29] = 1;cactus_sprite[0][25][30] = 1;cactus_sprite[0][25][31] = 1;cactus_sprite[0][25][32] = 1;cactus_sprite[0][25][33] = 1;cactus_sprite[0][25][34] = 1;cactus_sprite[0][25][35] = 1;cactus_sprite[0][25][36] = 1;cactus_sprite[0][25][37] = 1;cactus_sprite[0][25][38] = 1;cactus_sprite[0][25][39] = 1;cactus_sprite[0][25][40] = 1;cactus_sprite[0][25][41] = 1;cactus_sprite[0][25][42] = 1;cactus_sprite[0][25][43] = 1;cactus_sprite[0][25][44] = 1;cactus_sprite[0][25][45] = 1;cactus_sprite[0][25][46] = 1;cactus_sprite[0][25][47] = 1;cactus_sprite[0][25][48] = 1;cactus_sprite[0][25][49] = 1;cactus_sprite[0][25][50] = 1;cactus_sprite[0][25][51] = 1;cactus_sprite[0][25][52] = 1;cactus_sprite[0][25][53] = 1;cactus_sprite[0][25][54] = 1;cactus_sprite[0][25][55] = 1;cactus_sprite[0][25][56] = 1;cactus_sprite[0][25][57] = 1;cactus_sprite[0][25][58] = 1;cactus_sprite[0][25][59] = 1;cactus_sprite[0][25][60] = 1;cactus_sprite[0][25][61] = 1;cactus_sprite[0][25][62] = 1;cactus_sprite[0][25][63] = 1;cactus_sprite[0][25][64] = 1;cactus_sprite[0][25][65] = 1;cactus_sprite[0][25][66] = 1;cactus_sprite[0][25][67] = 1;cactus_sprite[0][25][68] = 1;cactus_sprite[0][25][69] = 1;cactus_sprite[0][25][70] = 1;cactus_sprite[0][25][71] = 1;cactus_sprite[0][25][72] = 1;cactus_sprite[0][25][73] = 1;cactus_sprite[0][25][74] = 1;cactus_sprite[0][25][75] = 1;cactus_sprite[0][25][76] = 1;cactus_sprite[0][25][77] = 1;cactus_sprite[0][25][78] = 1;cactus_sprite[0][25][79] = 1;cactus_sprite[0][25][80] = 1;cactus_sprite[0][25][81] = 1;cactus_sprite[0][25][82] = 1;cactus_sprite[0][25][83] = 1;cactus_sprite[0][25][84] = 1;cactus_sprite[0][25][85] = 1;cactus_sprite[0][25][86] = 1;cactus_sprite[0][25][87] = 1;cactus_sprite[0][25][88] = 1;cactus_sprite[0][25][89] = 1;cactus_sprite[0][25][90] = 1;cactus_sprite[0][25][91] = 1;cactus_sprite[0][25][92] = 1;cactus_sprite[0][25][93] = 1;cactus_sprite[0][25][94] = 1;cactus_sprite[0][25][95] = 1;cactus_sprite[0][25][96] = 1;cactus_sprite[0][25][97] = 1;cactus_sprite[0][25][98] = 1;cactus_sprite[0][25][99] = 1;cactus_sprite[0][26][8] = 1;cactus_sprite[0][26][9] = 1;cactus_sprite[0][26][10] = 1;cactus_sprite[0][26][11] = 1;cactus_sprite[0][26][12] = 1;cactus_sprite[0][26][13] = 1;cactus_sprite[0][26][14] = 1;cactus_sprite[0][26][15] = 1;cactus_sprite[0][26][16] = 1;cactus_sprite[0][26][17] = 1;cactus_sprite[0][26][18] = 1;cactus_sprite[0][26][19] = 1;cactus_sprite[0][26][20] = 1;cactus_sprite[0][26][21] = 1;cactus_sprite[0][26][22] = 1;cactus_sprite[0][26][23] = 1;cactus_sprite[0][26][24] = 1;cactus_sprite[0][26][25] = 1;cactus_sprite[0][26][26] = 1;cactus_sprite[0][26][27] = 1;cactus_sprite[0][26][28] = 1;cactus_sprite[0][26][29] = 1;cactus_sprite[0][26][30] = 1;cactus_sprite[0][26][31] = 1;cactus_sprite[0][26][32] = 1;cactus_sprite[0][26][33] = 1;cactus_sprite[0][26][34] = 1;cactus_sprite[0][26][35] = 1;cactus_sprite[0][26][36] = 1;cactus_sprite[0][26][37] = 1;cactus_sprite[0][26][38] = 1;cactus_sprite[0][26][39] = 1;cactus_sprite[0][26][40] = 1;cactus_sprite[0][26][41] = 1;cactus_sprite[0][26][42] = 1;cactus_sprite[0][26][43] = 1;cactus_sprite[0][26][44] = 1;cactus_sprite[0][26][45] = 1;cactus_sprite[0][26][46] = 1;cactus_sprite[0][26][47] = 1;cactus_sprite[0][26][48] = 1;cactus_sprite[0][26][49] = 1;cactus_sprite[0][26][50] = 1;cactus_sprite[0][26][51] = 1;cactus_sprite[0][26][52] = 1;cactus_sprite[0][26][53] = 1;cactus_sprite[0][26][54] = 1;cactus_sprite[0][26][55] = 1;cactus_sprite[0][26][56] = 1;cactus_sprite[0][26][57] = 1;cactus_sprite[0][26][58] = 1;cactus_sprite[0][26][59] = 1;cactus_sprite[0][26][60] = 1;cactus_sprite[0][26][61] = 1;cactus_sprite[0][26][62] = 1;cactus_sprite[0][26][63] = 1;cactus_sprite[0][26][64] = 1;cactus_sprite[0][26][65] = 1;cactus_sprite[0][26][66] = 1;cactus_sprite[0][26][67] = 1;cactus_sprite[0][26][68] = 1;cactus_sprite[0][26][69] = 1;cactus_sprite[0][26][70] = 1;cactus_sprite[0][26][71] = 1;cactus_sprite[0][26][72] = 1;cactus_sprite[0][26][73] = 1;cactus_sprite[0][26][74] = 1;cactus_sprite[0][26][75] = 1;cactus_sprite[0][26][76] = 1;cactus_sprite[0][26][77] = 1;cactus_sprite[0][26][78] = 1;cactus_sprite[0][26][79] = 1;cactus_sprite[0][26][80] = 1;cactus_sprite[0][26][81] = 1;cactus_sprite[0][26][82] = 1;cactus_sprite[0][26][83] = 1;cactus_sprite[0][26][84] = 1;cactus_sprite[0][26][85] = 1;cactus_sprite[0][26][86] = 1;cactus_sprite[0][26][87] = 1;cactus_sprite[0][26][88] = 1;cactus_sprite[0][26][89] = 1;cactus_sprite[0][26][90] = 1;cactus_sprite[0][26][91] = 1;cactus_sprite[0][26][92] = 1;cactus_sprite[0][26][93] = 1;cactus_sprite[0][26][94] = 1;cactus_sprite[0][26][95] = 1;cactus_sprite[0][26][96] = 1;cactus_sprite[0][26][97] = 1;cactus_sprite[0][26][98] = 1;cactus_sprite[0][26][99] = 1;cactus_sprite[0][27][8] = 1;cactus_sprite[0][27][9] = 1;cactus_sprite[0][27][10] = 1;cactus_sprite[0][27][11] = 1;cactus_sprite[0][27][12] = 1;cactus_sprite[0][27][13] = 1;cactus_sprite[0][27][14] = 1;cactus_sprite[0][27][15] = 1;cactus_sprite[0][27][16] = 1;cactus_sprite[0][27][17] = 1;cactus_sprite[0][27][18] = 1;cactus_sprite[0][27][19] = 1;cactus_sprite[0][27][20] = 1;cactus_sprite[0][27][21] = 1;cactus_sprite[0][27][22] = 1;cactus_sprite[0][27][23] = 1;cactus_sprite[0][27][24] = 1;cactus_sprite[0][27][25] = 1;cactus_sprite[0][27][26] = 1;cactus_sprite[0][27][27] = 1;cactus_sprite[0][27][28] = 1;cactus_sprite[0][27][29] = 1;cactus_sprite[0][27][30] = 1;cactus_sprite[0][27][31] = 1;cactus_sprite[0][27][32] = 1;cactus_sprite[0][27][33] = 1;cactus_sprite[0][27][34] = 1;cactus_sprite[0][27][35] = 1;cactus_sprite[0][27][36] = 1;cactus_sprite[0][27][37] = 1;cactus_sprite[0][27][38] = 1;cactus_sprite[0][27][39] = 1;cactus_sprite[0][27][40] = 1;cactus_sprite[0][27][41] = 1;cactus_sprite[0][27][42] = 1;cactus_sprite[0][27][43] = 1;cactus_sprite[0][27][44] = 1;cactus_sprite[0][27][45] = 1;cactus_sprite[0][27][46] = 1;cactus_sprite[0][27][47] = 1;cactus_sprite[0][27][48] = 1;cactus_sprite[0][27][49] = 1;cactus_sprite[0][27][50] = 1;cactus_sprite[0][27][51] = 1;cactus_sprite[0][27][52] = 1;cactus_sprite[0][27][53] = 1;cactus_sprite[0][27][54] = 1;cactus_sprite[0][27][55] = 1;cactus_sprite[0][27][56] = 1;cactus_sprite[0][27][57] = 1;cactus_sprite[0][27][58] = 1;cactus_sprite[0][27][59] = 1;cactus_sprite[0][27][60] = 1;cactus_sprite[0][27][61] = 1;cactus_sprite[0][27][62] = 1;cactus_sprite[0][27][63] = 1;cactus_sprite[0][27][64] = 1;cactus_sprite[0][27][65] = 1;cactus_sprite[0][27][66] = 1;cactus_sprite[0][27][67] = 1;cactus_sprite[0][27][68] = 1;cactus_sprite[0][27][69] = 1;cactus_sprite[0][27][70] = 1;cactus_sprite[0][27][71] = 1;cactus_sprite[0][27][72] = 1;cactus_sprite[0][27][73] = 1;cactus_sprite[0][27][74] = 1;cactus_sprite[0][27][75] = 1;cactus_sprite[0][27][76] = 1;cactus_sprite[0][27][77] = 1;cactus_sprite[0][27][78] = 1;cactus_sprite[0][27][79] = 1;cactus_sprite[0][27][80] = 1;cactus_sprite[0][27][81] = 1;cactus_sprite[0][27][82] = 1;cactus_sprite[0][27][83] = 1;cactus_sprite[0][27][84] = 1;cactus_sprite[0][27][85] = 1;cactus_sprite[0][27][86] = 1;cactus_sprite[0][27][87] = 1;cactus_sprite[0][27][88] = 1;cactus_sprite[0][27][89] = 1;cactus_sprite[0][27][90] = 1;cactus_sprite[0][27][91] = 1;cactus_sprite[0][27][92] = 1;cactus_sprite[0][27][93] = 1;cactus_sprite[0][27][94] = 1;cactus_sprite[0][27][95] = 1;cactus_sprite[0][27][96] = 1;cactus_sprite[0][27][97] = 1;cactus_sprite[0][27][98] = 1;cactus_sprite[0][27][99] = 1;cactus_sprite[0][28][8] = 1;cactus_sprite[0][28][9] = 1;cactus_sprite[0][28][10] = 1;cactus_sprite[0][28][11] = 1;cactus_sprite[0][28][12] = 1;cactus_sprite[0][28][13] = 1;cactus_sprite[0][28][14] = 1;cactus_sprite[0][28][15] = 1;cactus_sprite[0][28][16] = 1;cactus_sprite[0][28][17] = 1;cactus_sprite[0][28][18] = 1;cactus_sprite[0][28][19] = 1;cactus_sprite[0][28][20] = 1;cactus_sprite[0][28][21] = 1;cactus_sprite[0][28][22] = 1;cactus_sprite[0][28][23] = 1;cactus_sprite[0][28][24] = 1;cactus_sprite[0][28][25] = 1;cactus_sprite[0][28][26] = 1;cactus_sprite[0][28][27] = 1;cactus_sprite[0][28][28] = 1;cactus_sprite[0][28][29] = 1;cactus_sprite[0][28][30] = 1;cactus_sprite[0][28][31] = 1;cactus_sprite[0][28][32] = 1;cactus_sprite[0][28][33] = 1;cactus_sprite[0][28][34] = 1;cactus_sprite[0][28][35] = 1;cactus_sprite[0][28][36] = 1;cactus_sprite[0][28][37] = 1;cactus_sprite[0][28][38] = 1;cactus_sprite[0][28][39] = 1;cactus_sprite[0][28][40] = 1;cactus_sprite[0][28][41] = 1;cactus_sprite[0][28][42] = 1;cactus_sprite[0][28][43] = 1;cactus_sprite[0][28][44] = 1;cactus_sprite[0][28][45] = 1;cactus_sprite[0][28][46] = 1;cactus_sprite[0][28][47] = 1;cactus_sprite[0][28][48] = 1;cactus_sprite[0][28][49] = 1;cactus_sprite[0][28][50] = 1;cactus_sprite[0][28][51] = 1;cactus_sprite[0][28][52] = 1;cactus_sprite[0][28][53] = 1;cactus_sprite[0][28][54] = 1;cactus_sprite[0][28][55] = 1;cactus_sprite[0][28][56] = 1;cactus_sprite[0][28][57] = 1;cactus_sprite[0][28][58] = 1;cactus_sprite[0][28][59] = 1;cactus_sprite[0][28][60] = 1;cactus_sprite[0][28][61] = 1;cactus_sprite[0][28][62] = 1;cactus_sprite[0][28][63] = 1;cactus_sprite[0][28][64] = 1;cactus_sprite[0][28][65] = 1;cactus_sprite[0][28][66] = 1;cactus_sprite[0][28][67] = 1;cactus_sprite[0][28][68] = 1;cactus_sprite[0][28][69] = 1;cactus_sprite[0][28][70] = 1;cactus_sprite[0][28][71] = 1;cactus_sprite[0][28][72] = 1;cactus_sprite[0][28][73] = 1;cactus_sprite[0][28][74] = 1;cactus_sprite[0][28][75] = 1;cactus_sprite[0][28][76] = 1;cactus_sprite[0][28][77] = 1;cactus_sprite[0][28][78] = 1;cactus_sprite[0][28][79] = 1;cactus_sprite[0][28][80] = 1;cactus_sprite[0][28][81] = 1;cactus_sprite[0][28][82] = 1;cactus_sprite[0][28][83] = 1;cactus_sprite[0][28][84] = 1;cactus_sprite[0][28][85] = 1;cactus_sprite[0][28][86] = 1;cactus_sprite[0][28][87] = 1;cactus_sprite[0][28][88] = 1;cactus_sprite[0][28][89] = 1;cactus_sprite[0][28][90] = 1;cactus_sprite[0][28][91] = 1;cactus_sprite[0][28][92] = 1;cactus_sprite[0][28][93] = 1;cactus_sprite[0][28][94] = 1;cactus_sprite[0][28][95] = 1;cactus_sprite[0][28][96] = 1;cactus_sprite[0][28][97] = 1;cactus_sprite[0][28][98] = 1;cactus_sprite[0][28][99] = 1;cactus_sprite[0][29][8] = 1;cactus_sprite[0][29][9] = 1;cactus_sprite[0][29][10] = 1;cactus_sprite[0][29][11] = 1;cactus_sprite[0][29][12] = 1;cactus_sprite[0][29][13] = 1;cactus_sprite[0][29][14] = 1;cactus_sprite[0][29][15] = 1;cactus_sprite[0][29][16] = 1;cactus_sprite[0][29][17] = 1;cactus_sprite[0][29][18] = 1;cactus_sprite[0][29][19] = 1;cactus_sprite[0][29][20] = 1;cactus_sprite[0][29][21] = 1;cactus_sprite[0][29][22] = 1;cactus_sprite[0][29][23] = 1;cactus_sprite[0][29][24] = 1;cactus_sprite[0][29][25] = 1;cactus_sprite[0][29][26] = 1;cactus_sprite[0][29][27] = 1;cactus_sprite[0][29][28] = 1;cactus_sprite[0][29][29] = 1;cactus_sprite[0][29][30] = 1;cactus_sprite[0][29][31] = 1;cactus_sprite[0][29][32] = 1;cactus_sprite[0][29][33] = 1;cactus_sprite[0][29][34] = 1;cactus_sprite[0][29][35] = 1;cactus_sprite[0][29][36] = 1;cactus_sprite[0][29][37] = 1;cactus_sprite[0][29][38] = 1;cactus_sprite[0][29][39] = 1;cactus_sprite[0][29][40] = 1;cactus_sprite[0][29][41] = 1;cactus_sprite[0][29][42] = 1;cactus_sprite[0][29][43] = 1;cactus_sprite[0][29][44] = 1;cactus_sprite[0][29][45] = 1;cactus_sprite[0][29][46] = 1;cactus_sprite[0][29][47] = 1;cactus_sprite[0][29][48] = 1;cactus_sprite[0][29][49] = 1;cactus_sprite[0][29][50] = 1;cactus_sprite[0][29][51] = 1;cactus_sprite[0][29][52] = 1;cactus_sprite[0][29][53] = 1;cactus_sprite[0][29][54] = 1;cactus_sprite[0][29][55] = 1;cactus_sprite[0][29][56] = 1;cactus_sprite[0][29][57] = 1;cactus_sprite[0][29][58] = 1;cactus_sprite[0][29][59] = 1;cactus_sprite[0][29][60] = 1;cactus_sprite[0][29][61] = 1;cactus_sprite[0][29][62] = 1;cactus_sprite[0][29][63] = 1;cactus_sprite[0][29][64] = 1;cactus_sprite[0][29][65] = 1;cactus_sprite[0][29][66] = 1;cactus_sprite[0][29][67] = 1;cactus_sprite[0][29][68] = 1;cactus_sprite[0][29][69] = 1;cactus_sprite[0][29][70] = 1;cactus_sprite[0][29][71] = 1;cactus_sprite[0][29][72] = 1;cactus_sprite[0][29][73] = 1;cactus_sprite[0][29][74] = 1;cactus_sprite[0][29][75] = 1;cactus_sprite[0][29][76] = 1;cactus_sprite[0][29][77] = 1;cactus_sprite[0][29][78] = 1;cactus_sprite[0][29][79] = 1;cactus_sprite[0][29][80] = 1;cactus_sprite[0][29][81] = 1;cactus_sprite[0][29][82] = 1;cactus_sprite[0][29][83] = 1;cactus_sprite[0][29][84] = 1;cactus_sprite[0][29][85] = 1;cactus_sprite[0][29][86] = 1;cactus_sprite[0][29][87] = 1;cactus_sprite[0][29][88] = 1;cactus_sprite[0][29][89] = 1;cactus_sprite[0][29][90] = 1;cactus_sprite[0][29][91] = 1;cactus_sprite[0][29][92] = 1;cactus_sprite[0][29][93] = 1;cactus_sprite[0][29][94] = 1;cactus_sprite[0][29][95] = 1;cactus_sprite[0][29][96] = 1;cactus_sprite[0][29][97] = 1;cactus_sprite[0][29][98] = 1;cactus_sprite[0][29][99] = 1;cactus_sprite[0][30][10] = 1;cactus_sprite[0][30][11] = 1;cactus_sprite[0][30][12] = 1;cactus_sprite[0][30][13] = 1;cactus_sprite[0][30][14] = 1;cactus_sprite[0][30][15] = 1;cactus_sprite[0][30][16] = 1;cactus_sprite[0][30][17] = 1;cactus_sprite[0][30][18] = 1;cactus_sprite[0][30][19] = 1;cactus_sprite[0][30][20] = 1;cactus_sprite[0][30][21] = 1;cactus_sprite[0][30][22] = 1;cactus_sprite[0][30][23] = 1;cactus_sprite[0][30][24] = 1;cactus_sprite[0][30][25] = 1;cactus_sprite[0][30][26] = 1;cactus_sprite[0][30][27] = 1;cactus_sprite[0][30][28] = 1;cactus_sprite[0][30][29] = 1;cactus_sprite[0][30][30] = 1;cactus_sprite[0][30][31] = 1;cactus_sprite[0][30][32] = 1;cactus_sprite[0][30][33] = 1;cactus_sprite[0][30][34] = 1;cactus_sprite[0][30][35] = 1;cactus_sprite[0][30][36] = 1;cactus_sprite[0][30][37] = 1;cactus_sprite[0][30][38] = 1;cactus_sprite[0][30][39] = 1;cactus_sprite[0][30][40] = 1;cactus_sprite[0][30][41] = 1;cactus_sprite[0][30][42] = 1;cactus_sprite[0][30][43] = 1;cactus_sprite[0][30][44] = 1;cactus_sprite[0][30][45] = 1;cactus_sprite[0][30][46] = 1;cactus_sprite[0][30][47] = 1;cactus_sprite[0][30][48] = 1;cactus_sprite[0][30][49] = 1;cactus_sprite[0][30][50] = 1;cactus_sprite[0][30][51] = 1;cactus_sprite[0][30][52] = 1;cactus_sprite[0][30][53] = 1;cactus_sprite[0][30][54] = 1;cactus_sprite[0][30][55] = 1;cactus_sprite[0][30][56] = 1;cactus_sprite[0][30][57] = 1;cactus_sprite[0][30][58] = 1;cactus_sprite[0][30][59] = 1;cactus_sprite[0][30][60] = 1;cactus_sprite[0][30][61] = 1;cactus_sprite[0][30][62] = 1;cactus_sprite[0][30][63] = 1;cactus_sprite[0][30][64] = 1;cactus_sprite[0][30][65] = 1;cactus_sprite[0][30][66] = 1;cactus_sprite[0][30][67] = 1;cactus_sprite[0][30][68] = 1;cactus_sprite[0][30][69] = 1;cactus_sprite[0][30][70] = 1;cactus_sprite[0][30][71] = 1;cactus_sprite[0][30][72] = 1;cactus_sprite[0][30][73] = 1;cactus_sprite[0][30][74] = 1;cactus_sprite[0][30][75] = 1;cactus_sprite[0][30][76] = 1;cactus_sprite[0][30][77] = 1;cactus_sprite[0][30][78] = 1;cactus_sprite[0][30][79] = 1;cactus_sprite[0][30][80] = 1;cactus_sprite[0][30][81] = 1;cactus_sprite[0][30][82] = 1;cactus_sprite[0][30][83] = 1;cactus_sprite[0][30][84] = 1;cactus_sprite[0][30][85] = 1;cactus_sprite[0][30][86] = 1;cactus_sprite[0][30][87] = 1;cactus_sprite[0][30][88] = 1;cactus_sprite[0][30][89] = 1;cactus_sprite[0][30][90] = 1;cactus_sprite[0][30][91] = 1;cactus_sprite[0][30][92] = 1;cactus_sprite[0][30][93] = 1;cactus_sprite[0][30][94] = 1;cactus_sprite[0][30][95] = 1;cactus_sprite[0][30][96] = 1;cactus_sprite[0][30][97] = 1;cactus_sprite[0][30][98] = 1;cactus_sprite[0][30][99] = 1;cactus_sprite[0][31][10] = 1;cactus_sprite[0][31][11] = 1;cactus_sprite[0][31][12] = 1;cactus_sprite[0][31][13] = 1;cactus_sprite[0][31][14] = 1;cactus_sprite[0][31][15] = 1;cactus_sprite[0][31][16] = 1;cactus_sprite[0][31][17] = 1;cactus_sprite[0][31][18] = 1;cactus_sprite[0][31][19] = 1;cactus_sprite[0][31][20] = 1;cactus_sprite[0][31][21] = 1;cactus_sprite[0][31][22] = 1;cactus_sprite[0][31][23] = 1;cactus_sprite[0][31][24] = 1;cactus_sprite[0][31][25] = 1;cactus_sprite[0][31][26] = 1;cactus_sprite[0][31][27] = 1;cactus_sprite[0][31][28] = 1;cactus_sprite[0][31][29] = 1;cactus_sprite[0][31][30] = 1;cactus_sprite[0][31][31] = 1;cactus_sprite[0][31][32] = 1;cactus_sprite[0][31][33] = 1;cactus_sprite[0][31][34] = 1;cactus_sprite[0][31][35] = 1;cactus_sprite[0][31][36] = 1;cactus_sprite[0][31][37] = 1;cactus_sprite[0][31][38] = 1;cactus_sprite[0][31][39] = 1;cactus_sprite[0][31][40] = 1;cactus_sprite[0][31][41] = 1;cactus_sprite[0][31][42] = 1;cactus_sprite[0][31][43] = 1;cactus_sprite[0][31][44] = 1;cactus_sprite[0][31][45] = 1;cactus_sprite[0][31][46] = 1;cactus_sprite[0][31][47] = 1;cactus_sprite[0][31][48] = 1;cactus_sprite[0][31][49] = 1;cactus_sprite[0][31][50] = 1;cactus_sprite[0][31][51] = 1;cactus_sprite[0][31][52] = 1;cactus_sprite[0][31][53] = 1;cactus_sprite[0][31][54] = 1;cactus_sprite[0][31][55] = 1;cactus_sprite[0][31][56] = 1;cactus_sprite[0][31][57] = 1;cactus_sprite[0][31][58] = 1;cactus_sprite[0][31][59] = 1;cactus_sprite[0][31][60] = 1;cactus_sprite[0][31][61] = 1;cactus_sprite[0][31][62] = 1;cactus_sprite[0][31][63] = 1;cactus_sprite[0][31][64] = 1;cactus_sprite[0][31][65] = 1;cactus_sprite[0][31][66] = 1;cactus_sprite[0][31][67] = 1;cactus_sprite[0][31][68] = 1;cactus_sprite[0][31][69] = 1;cactus_sprite[0][31][70] = 1;cactus_sprite[0][31][71] = 1;cactus_sprite[0][31][72] = 1;cactus_sprite[0][31][73] = 1;cactus_sprite[0][31][74] = 1;cactus_sprite[0][31][75] = 1;cactus_sprite[0][31][76] = 1;cactus_sprite[0][31][77] = 1;cactus_sprite[0][31][78] = 1;cactus_sprite[0][31][79] = 1;cactus_sprite[0][31][80] = 1;cactus_sprite[0][31][81] = 1;cactus_sprite[0][31][82] = 1;cactus_sprite[0][31][83] = 1;cactus_sprite[0][31][84] = 1;cactus_sprite[0][31][85] = 1;cactus_sprite[0][31][86] = 1;cactus_sprite[0][31][87] = 1;cactus_sprite[0][31][88] = 1;cactus_sprite[0][31][89] = 1;cactus_sprite[0][31][90] = 1;cactus_sprite[0][31][91] = 1;cactus_sprite[0][31][92] = 1;cactus_sprite[0][31][93] = 1;cactus_sprite[0][31][94] = 1;cactus_sprite[0][31][95] = 1;cactus_sprite[0][31][96] = 1;cactus_sprite[0][31][97] = 1;cactus_sprite[0][31][98] = 1;cactus_sprite[0][31][99] = 1;cactus_sprite[0][32][60] = 1;cactus_sprite[0][32][61] = 1;cactus_sprite[0][32][62] = 1;cactus_sprite[0][32][63] = 1;cactus_sprite[0][32][64] = 1;cactus_sprite[0][32][65] = 1;cactus_sprite[0][32][66] = 1;cactus_sprite[0][32][67] = 1;cactus_sprite[0][33][60] = 1;cactus_sprite[0][33][61] = 1;cactus_sprite[0][33][62] = 1;cactus_sprite[0][33][63] = 1;cactus_sprite[0][33][64] = 1;cactus_sprite[0][33][65] = 1;cactus_sprite[0][33][66] = 1;cactus_sprite[0][33][67] = 1;cactus_sprite[0][34][60] = 1;cactus_sprite[0][34][61] = 1;cactus_sprite[0][34][62] = 1;cactus_sprite[0][34][63] = 1;cactus_sprite[0][34][64] = 1;cactus_sprite[0][34][65] = 1;cactus_sprite[0][34][66] = 1;cactus_sprite[0][34][67] = 1;cactus_sprite[0][35][60] = 1;cactus_sprite[0][35][61] = 1;cactus_sprite[0][35][62] = 1;cactus_sprite[0][35][63] = 1;cactus_sprite[0][35][64] = 1;cactus_sprite[0][35][65] = 1;cactus_sprite[0][35][66] = 1;cactus_sprite[0][35][67] = 1;cactus_sprite[0][36][60] = 1;cactus_sprite[0][36][61] = 1;cactus_sprite[0][36][62] = 1;cactus_sprite[0][36][63] = 1;cactus_sprite[0][36][64] = 1;cactus_sprite[0][36][65] = 1;cactus_sprite[0][36][66] = 1;cactus_sprite[0][36][67] = 1;cactus_sprite[0][37][60] = 1;cactus_sprite[0][37][61] = 1;cactus_sprite[0][37][62] = 1;cactus_sprite[0][37][63] = 1;cactus_sprite[0][37][64] = 1;cactus_sprite[0][37][65] = 1;cactus_sprite[0][37][66] = 1;cactus_sprite[0][37][67] = 1;cactus_sprite[0][38][30] = 1;cactus_sprite[0][38][31] = 1;cactus_sprite[0][38][32] = 1;cactus_sprite[0][38][33] = 1;cactus_sprite[0][38][34] = 1;cactus_sprite[0][38][35] = 1;cactus_sprite[0][38][36] = 1;cactus_sprite[0][38][37] = 1;cactus_sprite[0][38][38] = 1;cactus_sprite[0][38][39] = 1;cactus_sprite[0][38][40] = 1;cactus_sprite[0][38][41] = 1;cactus_sprite[0][38][42] = 1;cactus_sprite[0][38][43] = 1;cactus_sprite[0][38][44] = 1;cactus_sprite[0][38][45] = 1;cactus_sprite[0][38][46] = 1;cactus_sprite[0][38][47] = 1;cactus_sprite[0][38][48] = 1;cactus_sprite[0][38][49] = 1;cactus_sprite[0][38][50] = 1;cactus_sprite[0][38][51] = 1;cactus_sprite[0][38][52] = 1;cactus_sprite[0][38][53] = 1;cactus_sprite[0][38][54] = 1;cactus_sprite[0][38][55] = 1;cactus_sprite[0][38][56] = 1;cactus_sprite[0][38][57] = 1;cactus_sprite[0][38][58] = 1;cactus_sprite[0][38][59] = 1;cactus_sprite[0][38][60] = 1;cactus_sprite[0][38][61] = 1;cactus_sprite[0][38][62] = 1;cactus_sprite[0][38][63] = 1;cactus_sprite[0][38][64] = 1;cactus_sprite[0][38][65] = 1;cactus_sprite[0][38][66] = 1;cactus_sprite[0][38][67] = 1;cactus_sprite[0][39][30] = 1;cactus_sprite[0][39][31] = 1;cactus_sprite[0][39][32] = 1;cactus_sprite[0][39][33] = 1;cactus_sprite[0][39][34] = 1;cactus_sprite[0][39][35] = 1;cactus_sprite[0][39][36] = 1;cactus_sprite[0][39][37] = 1;cactus_sprite[0][39][38] = 1;cactus_sprite[0][39][39] = 1;cactus_sprite[0][39][40] = 1;cactus_sprite[0][39][41] = 1;cactus_sprite[0][39][42] = 1;cactus_sprite[0][39][43] = 1;cactus_sprite[0][39][44] = 1;cactus_sprite[0][39][45] = 1;cactus_sprite[0][39][46] = 1;cactus_sprite[0][39][47] = 1;cactus_sprite[0][39][48] = 1;cactus_sprite[0][39][49] = 1;cactus_sprite[0][39][50] = 1;cactus_sprite[0][39][51] = 1;cactus_sprite[0][39][52] = 1;cactus_sprite[0][39][53] = 1;cactus_sprite[0][39][54] = 1;cactus_sprite[0][39][55] = 1;cactus_sprite[0][39][56] = 1;cactus_sprite[0][39][57] = 1;cactus_sprite[0][39][58] = 1;cactus_sprite[0][39][59] = 1;cactus_sprite[0][39][60] = 1;cactus_sprite[0][39][61] = 1;cactus_sprite[0][39][62] = 1;cactus_sprite[0][39][63] = 1;cactus_sprite[0][39][64] = 1;cactus_sprite[0][39][65] = 1;cactus_sprite[0][39][66] = 1;cactus_sprite[0][39][67] = 1;cactus_sprite[0][40][28] = 1;cactus_sprite[0][40][29] = 1;cactus_sprite[0][40][30] = 1;cactus_sprite[0][40][31] = 1;cactus_sprite[0][40][32] = 1;cactus_sprite[0][40][33] = 1;cactus_sprite[0][40][34] = 1;cactus_sprite[0][40][35] = 1;cactus_sprite[0][40][36] = 1;cactus_sprite[0][40][37] = 1;cactus_sprite[0][40][38] = 1;cactus_sprite[0][40][39] = 1;cactus_sprite[0][40][40] = 1;cactus_sprite[0][40][41] = 1;cactus_sprite[0][40][42] = 1;cactus_sprite[0][40][43] = 1;cactus_sprite[0][40][44] = 1;cactus_sprite[0][40][45] = 1;cactus_sprite[0][40][46] = 1;cactus_sprite[0][40][47] = 1;cactus_sprite[0][40][48] = 1;cactus_sprite[0][40][49] = 1;cactus_sprite[0][40][50] = 1;cactus_sprite[0][40][51] = 1;cactus_sprite[0][40][52] = 1;cactus_sprite[0][40][53] = 1;cactus_sprite[0][40][54] = 1;cactus_sprite[0][40][55] = 1;cactus_sprite[0][40][56] = 1;cactus_sprite[0][40][57] = 1;cactus_sprite[0][40][58] = 1;cactus_sprite[0][40][59] = 1;cactus_sprite[0][40][60] = 1;cactus_sprite[0][40][61] = 1;cactus_sprite[0][40][62] = 1;cactus_sprite[0][40][63] = 1;cactus_sprite[0][40][64] = 1;cactus_sprite[0][40][65] = 1;cactus_sprite[0][41][28] = 1;cactus_sprite[0][41][29] = 1;cactus_sprite[0][41][30] = 1;cactus_sprite[0][41][31] = 1;cactus_sprite[0][41][32] = 1;cactus_sprite[0][41][33] = 1;cactus_sprite[0][41][34] = 1;cactus_sprite[0][41][35] = 1;cactus_sprite[0][41][36] = 1;cactus_sprite[0][41][37] = 1;cactus_sprite[0][41][38] = 1;cactus_sprite[0][41][39] = 1;cactus_sprite[0][41][40] = 1;cactus_sprite[0][41][41] = 1;cactus_sprite[0][41][42] = 1;cactus_sprite[0][41][43] = 1;cactus_sprite[0][41][44] = 1;cactus_sprite[0][41][45] = 1;cactus_sprite[0][41][46] = 1;cactus_sprite[0][41][47] = 1;cactus_sprite[0][41][48] = 1;cactus_sprite[0][41][49] = 1;cactus_sprite[0][41][50] = 1;cactus_sprite[0][41][51] = 1;cactus_sprite[0][41][52] = 1;cactus_sprite[0][41][53] = 1;cactus_sprite[0][41][54] = 1;cactus_sprite[0][41][55] = 1;cactus_sprite[0][41][56] = 1;cactus_sprite[0][41][57] = 1;cactus_sprite[0][41][58] = 1;cactus_sprite[0][41][59] = 1;cactus_sprite[0][41][60] = 1;cactus_sprite[0][41][61] = 1;cactus_sprite[0][41][62] = 1;cactus_sprite[0][41][63] = 1;cactus_sprite[0][41][64] = 1;cactus_sprite[0][41][65] = 1;cactus_sprite[0][42][28] = 1;cactus_sprite[0][42][29] = 1;cactus_sprite[0][42][30] = 1;cactus_sprite[0][42][31] = 1;cactus_sprite[0][42][32] = 1;cactus_sprite[0][42][33] = 1;cactus_sprite[0][42][34] = 1;cactus_sprite[0][42][35] = 1;cactus_sprite[0][42][36] = 1;cactus_sprite[0][42][37] = 1;cactus_sprite[0][42][38] = 1;cactus_sprite[0][42][39] = 1;cactus_sprite[0][42][40] = 1;cactus_sprite[0][42][41] = 1;cactus_sprite[0][42][42] = 1;cactus_sprite[0][42][43] = 1;cactus_sprite[0][42][44] = 1;cactus_sprite[0][42][45] = 1;cactus_sprite[0][42][46] = 1;cactus_sprite[0][42][47] = 1;cactus_sprite[0][42][48] = 1;cactus_sprite[0][42][49] = 1;cactus_sprite[0][42][50] = 1;cactus_sprite[0][42][51] = 1;cactus_sprite[0][42][52] = 1;cactus_sprite[0][42][53] = 1;cactus_sprite[0][42][54] = 1;cactus_sprite[0][42][55] = 1;cactus_sprite[0][42][56] = 1;cactus_sprite[0][42][57] = 1;cactus_sprite[0][42][58] = 1;cactus_sprite[0][42][59] = 1;cactus_sprite[0][42][60] = 1;cactus_sprite[0][42][61] = 1;cactus_sprite[0][42][62] = 1;cactus_sprite[0][42][63] = 1;cactus_sprite[0][43][28] = 1;cactus_sprite[0][43][29] = 1;cactus_sprite[0][43][30] = 1;cactus_sprite[0][43][31] = 1;cactus_sprite[0][43][32] = 1;cactus_sprite[0][43][33] = 1;cactus_sprite[0][43][34] = 1;cactus_sprite[0][43][35] = 1;cactus_sprite[0][43][36] = 1;cactus_sprite[0][43][37] = 1;cactus_sprite[0][43][38] = 1;cactus_sprite[0][43][39] = 1;cactus_sprite[0][43][40] = 1;cactus_sprite[0][43][41] = 1;cactus_sprite[0][43][42] = 1;cactus_sprite[0][43][43] = 1;cactus_sprite[0][43][44] = 1;cactus_sprite[0][43][45] = 1;cactus_sprite[0][43][46] = 1;cactus_sprite[0][43][47] = 1;cactus_sprite[0][43][48] = 1;cactus_sprite[0][43][49] = 1;cactus_sprite[0][43][50] = 1;cactus_sprite[0][43][51] = 1;cactus_sprite[0][43][52] = 1;cactus_sprite[0][43][53] = 1;cactus_sprite[0][43][54] = 1;cactus_sprite[0][43][55] = 1;cactus_sprite[0][43][56] = 1;cactus_sprite[0][43][57] = 1;cactus_sprite[0][43][58] = 1;cactus_sprite[0][43][59] = 1;cactus_sprite[0][43][60] = 1;cactus_sprite[0][43][61] = 1;cactus_sprite[0][43][62] = 1;cactus_sprite[0][43][63] = 1;cactus_sprite[0][44][28] = 1;cactus_sprite[0][44][29] = 1;cactus_sprite[0][44][30] = 1;cactus_sprite[0][44][31] = 1;cactus_sprite[0][44][32] = 1;cactus_sprite[0][44][33] = 1;cactus_sprite[0][44][34] = 1;cactus_sprite[0][44][35] = 1;cactus_sprite[0][44][36] = 1;cactus_sprite[0][44][37] = 1;cactus_sprite[0][44][38] = 1;cactus_sprite[0][44][39] = 1;cactus_sprite[0][44][40] = 1;cactus_sprite[0][44][41] = 1;cactus_sprite[0][44][42] = 1;cactus_sprite[0][44][43] = 1;cactus_sprite[0][44][44] = 1;cactus_sprite[0][44][45] = 1;cactus_sprite[0][44][46] = 1;cactus_sprite[0][44][47] = 1;cactus_sprite[0][44][48] = 1;cactus_sprite[0][44][49] = 1;cactus_sprite[0][44][50] = 1;cactus_sprite[0][44][51] = 1;cactus_sprite[0][44][52] = 1;cactus_sprite[0][44][53] = 1;cactus_sprite[0][44][54] = 1;cactus_sprite[0][44][55] = 1;cactus_sprite[0][44][56] = 1;cactus_sprite[0][44][57] = 1;cactus_sprite[0][44][58] = 1;cactus_sprite[0][44][59] = 1;cactus_sprite[0][44][60] = 1;cactus_sprite[0][44][61] = 1;cactus_sprite[0][45][28] = 1;cactus_sprite[0][45][29] = 1;cactus_sprite[0][45][30] = 1;cactus_sprite[0][45][31] = 1;cactus_sprite[0][45][32] = 1;cactus_sprite[0][45][33] = 1;cactus_sprite[0][45][34] = 1;cactus_sprite[0][45][35] = 1;cactus_sprite[0][45][36] = 1;cactus_sprite[0][45][37] = 1;cactus_sprite[0][45][38] = 1;cactus_sprite[0][45][39] = 1;cactus_sprite[0][45][40] = 1;cactus_sprite[0][45][41] = 1;cactus_sprite[0][45][42] = 1;cactus_sprite[0][45][43] = 1;cactus_sprite[0][45][44] = 1;cactus_sprite[0][45][45] = 1;cactus_sprite[0][45][46] = 1;cactus_sprite[0][45][47] = 1;cactus_sprite[0][45][48] = 1;cactus_sprite[0][45][49] = 1;cactus_sprite[0][45][50] = 1;cactus_sprite[0][45][51] = 1;cactus_sprite[0][45][52] = 1;cactus_sprite[0][45][53] = 1;cactus_sprite[0][45][54] = 1;cactus_sprite[0][45][55] = 1;cactus_sprite[0][45][56] = 1;cactus_sprite[0][45][57] = 1;cactus_sprite[0][45][58] = 1;cactus_sprite[0][45][59] = 1;cactus_sprite[0][45][60] = 1;cactus_sprite[0][45][61] = 1;cactus_sprite[0][46][30] = 1;cactus_sprite[0][46][31] = 1;cactus_sprite[0][46][32] = 1;cactus_sprite[0][46][33] = 1;cactus_sprite[0][46][34] = 1;cactus_sprite[0][46][35] = 1;cactus_sprite[0][46][36] = 1;cactus_sprite[0][46][37] = 1;cactus_sprite[0][46][38] = 1;cactus_sprite[0][46][39] = 1;cactus_sprite[0][46][40] = 1;cactus_sprite[0][46][41] = 1;cactus_sprite[0][46][42] = 1;cactus_sprite[0][46][43] = 1;cactus_sprite[0][46][44] = 1;cactus_sprite[0][46][45] = 1;cactus_sprite[0][46][46] = 1;cactus_sprite[0][46][47] = 1;cactus_sprite[0][46][48] = 1;cactus_sprite[0][46][49] = 1;cactus_sprite[0][46][50] = 1;cactus_sprite[0][46][51] = 1;cactus_sprite[0][46][52] = 1;cactus_sprite[0][46][53] = 1;cactus_sprite[0][46][54] = 1;cactus_sprite[0][46][55] = 1;cactus_sprite[0][46][56] = 1;cactus_sprite[0][46][57] = 1;cactus_sprite[0][46][58] = 1;cactus_sprite[0][46][59] = 1;cactus_sprite[0][47][30] = 1;cactus_sprite[0][47][31] = 1;cactus_sprite[0][47][32] = 1;cactus_sprite[0][47][33] = 1;cactus_sprite[0][47][34] = 1;cactus_sprite[0][47][35] = 1;cactus_sprite[0][47][36] = 1;cactus_sprite[0][47][37] = 1;cactus_sprite[0][47][38] = 1;cactus_sprite[0][47][39] = 1;cactus_sprite[0][47][40] = 1;cactus_sprite[0][47][41] = 1;cactus_sprite[0][47][42] = 1;cactus_sprite[0][47][43] = 1;cactus_sprite[0][47][44] = 1;cactus_sprite[0][47][45] = 1;cactus_sprite[0][47][46] = 1;cactus_sprite[0][47][47] = 1;cactus_sprite[0][47][48] = 1;cactus_sprite[0][47][49] = 1;cactus_sprite[0][47][50] = 1;cactus_sprite[0][47][51] = 1;cactus_sprite[0][47][52] = 1;cactus_sprite[0][47][53] = 1;cactus_sprite[0][47][54] = 1;cactus_sprite[0][47][55] = 1;cactus_sprite[0][47][56] = 1;cactus_sprite[0][47][57] = 1;cactus_sprite[0][47][58] = 1;cactus_sprite[0][47][59] = 1;
	cactus_sprite[1][2][34] = 1;cactus_sprite[1][2][35] = 1;cactus_sprite[1][2][36] = 1;cactus_sprite[1][2][37] = 1;cactus_sprite[1][2][38] = 1;cactus_sprite[1][2][39] = 1;cactus_sprite[1][2][40] = 1;cactus_sprite[1][2][41] = 1;cactus_sprite[1][2][42] = 1;cactus_sprite[1][2][43] = 1;cactus_sprite[1][2][44] = 1;cactus_sprite[1][2][45] = 1;cactus_sprite[1][2][46] = 1;cactus_sprite[1][2][47] = 1;cactus_sprite[1][2][48] = 1;cactus_sprite[1][2][49] = 1;cactus_sprite[1][2][50] = 1;cactus_sprite[1][2][51] = 1;cactus_sprite[1][2][52] = 1;cactus_sprite[1][2][53] = 1;cactus_sprite[1][2][54] = 1;cactus_sprite[1][2][55] = 1;cactus_sprite[1][2][56] = 1;cactus_sprite[1][2][57] = 1;cactus_sprite[1][2][58] = 1;cactus_sprite[1][2][59] = 1;cactus_sprite[1][2][60] = 1;cactus_sprite[1][2][61] = 1;cactus_sprite[1][2][62] = 1;cactus_sprite[1][2][63] = 1;cactus_sprite[1][3][34] = 1;cactus_sprite[1][3][35] = 1;cactus_sprite[1][3][36] = 1;cactus_sprite[1][3][37] = 1;cactus_sprite[1][3][38] = 1;cactus_sprite[1][3][39] = 1;cactus_sprite[1][3][40] = 1;cactus_sprite[1][3][41] = 1;cactus_sprite[1][3][42] = 1;cactus_sprite[1][3][43] = 1;cactus_sprite[1][3][44] = 1;cactus_sprite[1][3][45] = 1;cactus_sprite[1][3][46] = 1;cactus_sprite[1][3][47] = 1;cactus_sprite[1][3][48] = 1;cactus_sprite[1][3][49] = 1;cactus_sprite[1][3][50] = 1;cactus_sprite[1][3][51] = 1;cactus_sprite[1][3][52] = 1;cactus_sprite[1][3][53] = 1;cactus_sprite[1][3][54] = 1;cactus_sprite[1][3][55] = 1;cactus_sprite[1][3][56] = 1;cactus_sprite[1][3][57] = 1;cactus_sprite[1][3][58] = 1;cactus_sprite[1][3][59] = 1;cactus_sprite[1][3][60] = 1;cactus_sprite[1][3][61] = 1;cactus_sprite[1][3][62] = 1;cactus_sprite[1][3][63] = 1;cactus_sprite[1][4][32] = 1;cactus_sprite[1][4][33] = 1;cactus_sprite[1][4][34] = 1;cactus_sprite[1][4][35] = 1;cactus_sprite[1][4][36] = 1;cactus_sprite[1][4][37] = 1;cactus_sprite[1][4][38] = 1;cactus_sprite[1][4][39] = 1;cactus_sprite[1][4][40] = 1;cactus_sprite[1][4][41] = 1;cactus_sprite[1][4][42] = 1;cactus_sprite[1][4][43] = 1;cactus_sprite[1][4][44] = 1;cactus_sprite[1][4][45] = 1;cactus_sprite[1][4][46] = 1;cactus_sprite[1][4][47] = 1;cactus_sprite[1][4][48] = 1;cactus_sprite[1][4][49] = 1;cactus_sprite[1][4][50] = 1;cactus_sprite[1][4][51] = 1;cactus_sprite[1][4][52] = 1;cactus_sprite[1][4][53] = 1;cactus_sprite[1][4][54] = 1;cactus_sprite[1][4][55] = 1;cactus_sprite[1][4][56] = 1;cactus_sprite[1][4][57] = 1;cactus_sprite[1][4][58] = 1;cactus_sprite[1][4][59] = 1;cactus_sprite[1][4][60] = 1;cactus_sprite[1][4][61] = 1;cactus_sprite[1][4][62] = 1;cactus_sprite[1][4][63] = 1;cactus_sprite[1][4][64] = 1;cactus_sprite[1][4][65] = 1;cactus_sprite[1][5][32] = 1;cactus_sprite[1][5][33] = 1;cactus_sprite[1][5][34] = 1;cactus_sprite[1][5][35] = 1;cactus_sprite[1][5][36] = 1;cactus_sprite[1][5][37] = 1;cactus_sprite[1][5][38] = 1;cactus_sprite[1][5][39] = 1;cactus_sprite[1][5][40] = 1;cactus_sprite[1][5][41] = 1;cactus_sprite[1][5][42] = 1;cactus_sprite[1][5][43] = 1;cactus_sprite[1][5][44] = 1;cactus_sprite[1][5][45] = 1;cactus_sprite[1][5][46] = 1;cactus_sprite[1][5][47] = 1;cactus_sprite[1][5][48] = 1;cactus_sprite[1][5][49] = 1;cactus_sprite[1][5][50] = 1;cactus_sprite[1][5][51] = 1;cactus_sprite[1][5][52] = 1;cactus_sprite[1][5][53] = 1;cactus_sprite[1][5][54] = 1;cactus_sprite[1][5][55] = 1;cactus_sprite[1][5][56] = 1;cactus_sprite[1][5][57] = 1;cactus_sprite[1][5][58] = 1;cactus_sprite[1][5][59] = 1;cactus_sprite[1][5][60] = 1;cactus_sprite[1][5][61] = 1;cactus_sprite[1][5][62] = 1;cactus_sprite[1][5][63] = 1;cactus_sprite[1][5][64] = 1;cactus_sprite[1][5][65] = 1;cactus_sprite[1][6][32] = 1;cactus_sprite[1][6][33] = 1;cactus_sprite[1][6][34] = 1;cactus_sprite[1][6][35] = 1;cactus_sprite[1][6][36] = 1;cactus_sprite[1][6][37] = 1;cactus_sprite[1][6][38] = 1;cactus_sprite[1][6][39] = 1;cactus_sprite[1][6][40] = 1;cactus_sprite[1][6][41] = 1;cactus_sprite[1][6][42] = 1;cactus_sprite[1][6][43] = 1;cactus_sprite[1][6][44] = 1;cactus_sprite[1][6][45] = 1;cactus_sprite[1][6][46] = 1;cactus_sprite[1][6][47] = 1;cactus_sprite[1][6][48] = 1;cactus_sprite[1][6][49] = 1;cactus_sprite[1][6][50] = 1;cactus_sprite[1][6][51] = 1;cactus_sprite[1][6][52] = 1;cactus_sprite[1][6][53] = 1;cactus_sprite[1][6][54] = 1;cactus_sprite[1][6][55] = 1;cactus_sprite[1][6][56] = 1;cactus_sprite[1][6][57] = 1;cactus_sprite[1][6][58] = 1;cactus_sprite[1][6][59] = 1;cactus_sprite[1][6][60] = 1;cactus_sprite[1][6][61] = 1;cactus_sprite[1][6][62] = 1;cactus_sprite[1][6][63] = 1;cactus_sprite[1][6][64] = 1;cactus_sprite[1][6][65] = 1;cactus_sprite[1][6][66] = 1;cactus_sprite[1][6][67] = 1;cactus_sprite[1][7][32] = 1;cactus_sprite[1][7][33] = 1;cactus_sprite[1][7][34] = 1;cactus_sprite[1][7][35] = 1;cactus_sprite[1][7][36] = 1;cactus_sprite[1][7][37] = 1;cactus_sprite[1][7][38] = 1;cactus_sprite[1][7][39] = 1;cactus_sprite[1][7][40] = 1;cactus_sprite[1][7][41] = 1;cactus_sprite[1][7][42] = 1;cactus_sprite[1][7][43] = 1;cactus_sprite[1][7][44] = 1;cactus_sprite[1][7][45] = 1;cactus_sprite[1][7][46] = 1;cactus_sprite[1][7][47] = 1;cactus_sprite[1][7][48] = 1;cactus_sprite[1][7][49] = 1;cactus_sprite[1][7][50] = 1;cactus_sprite[1][7][51] = 1;cactus_sprite[1][7][52] = 1;cactus_sprite[1][7][53] = 1;cactus_sprite[1][7][54] = 1;cactus_sprite[1][7][55] = 1;cactus_sprite[1][7][56] = 1;cactus_sprite[1][7][57] = 1;cactus_sprite[1][7][58] = 1;cactus_sprite[1][7][59] = 1;cactus_sprite[1][7][60] = 1;cactus_sprite[1][7][61] = 1;cactus_sprite[1][7][62] = 1;cactus_sprite[1][7][63] = 1;cactus_sprite[1][7][64] = 1;cactus_sprite[1][7][65] = 1;cactus_sprite[1][7][66] = 1;cactus_sprite[1][7][67] = 1;cactus_sprite[1][8][32] = 1;cactus_sprite[1][8][33] = 1;cactus_sprite[1][8][34] = 1;cactus_sprite[1][8][35] = 1;cactus_sprite[1][8][36] = 1;cactus_sprite[1][8][37] = 1;cactus_sprite[1][8][38] = 1;cactus_sprite[1][8][39] = 1;cactus_sprite[1][8][40] = 1;cactus_sprite[1][8][41] = 1;cactus_sprite[1][8][42] = 1;cactus_sprite[1][8][43] = 1;cactus_sprite[1][8][44] = 1;cactus_sprite[1][8][45] = 1;cactus_sprite[1][8][46] = 1;cactus_sprite[1][8][47] = 1;cactus_sprite[1][8][48] = 1;cactus_sprite[1][8][49] = 1;cactus_sprite[1][8][50] = 1;cactus_sprite[1][8][51] = 1;cactus_sprite[1][8][52] = 1;cactus_sprite[1][8][53] = 1;cactus_sprite[1][8][54] = 1;cactus_sprite[1][8][55] = 1;cactus_sprite[1][8][56] = 1;cactus_sprite[1][8][57] = 1;cactus_sprite[1][8][58] = 1;cactus_sprite[1][8][59] = 1;cactus_sprite[1][8][60] = 1;cactus_sprite[1][8][61] = 1;cactus_sprite[1][8][62] = 1;cactus_sprite[1][8][63] = 1;cactus_sprite[1][8][64] = 1;cactus_sprite[1][8][65] = 1;cactus_sprite[1][8][66] = 1;cactus_sprite[1][8][67] = 1;cactus_sprite[1][8][68] = 1;cactus_sprite[1][8][69] = 1;cactus_sprite[1][9][32] = 1;cactus_sprite[1][9][33] = 1;cactus_sprite[1][9][34] = 1;cactus_sprite[1][9][35] = 1;cactus_sprite[1][9][36] = 1;cactus_sprite[1][9][37] = 1;cactus_sprite[1][9][38] = 1;cactus_sprite[1][9][39] = 1;cactus_sprite[1][9][40] = 1;cactus_sprite[1][9][41] = 1;cactus_sprite[1][9][42] = 1;cactus_sprite[1][9][43] = 1;cactus_sprite[1][9][44] = 1;cactus_sprite[1][9][45] = 1;cactus_sprite[1][9][46] = 1;cactus_sprite[1][9][47] = 1;cactus_sprite[1][9][48] = 1;cactus_sprite[1][9][49] = 1;cactus_sprite[1][9][50] = 1;cactus_sprite[1][9][51] = 1;cactus_sprite[1][9][52] = 1;cactus_sprite[1][9][53] = 1;cactus_sprite[1][9][54] = 1;cactus_sprite[1][9][55] = 1;cactus_sprite[1][9][56] = 1;cactus_sprite[1][9][57] = 1;cactus_sprite[1][9][58] = 1;cactus_sprite[1][9][59] = 1;cactus_sprite[1][9][60] = 1;cactus_sprite[1][9][61] = 1;cactus_sprite[1][9][62] = 1;cactus_sprite[1][9][63] = 1;cactus_sprite[1][9][64] = 1;cactus_sprite[1][9][65] = 1;cactus_sprite[1][9][66] = 1;cactus_sprite[1][9][67] = 1;cactus_sprite[1][9][68] = 1;cactus_sprite[1][9][69] = 1;cactus_sprite[1][10][34] = 1;cactus_sprite[1][10][35] = 1;cactus_sprite[1][10][36] = 1;cactus_sprite[1][10][37] = 1;cactus_sprite[1][10][38] = 1;cactus_sprite[1][10][39] = 1;cactus_sprite[1][10][40] = 1;cactus_sprite[1][10][41] = 1;cactus_sprite[1][10][42] = 1;cactus_sprite[1][10][43] = 1;cactus_sprite[1][10][44] = 1;cactus_sprite[1][10][45] = 1;cactus_sprite[1][10][46] = 1;cactus_sprite[1][10][47] = 1;cactus_sprite[1][10][48] = 1;cactus_sprite[1][10][49] = 1;cactus_sprite[1][10][50] = 1;cactus_sprite[1][10][51] = 1;cactus_sprite[1][10][52] = 1;cactus_sprite[1][10][53] = 1;cactus_sprite[1][10][54] = 1;cactus_sprite[1][10][55] = 1;cactus_sprite[1][10][56] = 1;cactus_sprite[1][10][57] = 1;cactus_sprite[1][10][58] = 1;cactus_sprite[1][10][59] = 1;cactus_sprite[1][10][60] = 1;cactus_sprite[1][10][61] = 1;cactus_sprite[1][10][62] = 1;cactus_sprite[1][10][63] = 1;cactus_sprite[1][10][64] = 1;cactus_sprite[1][10][65] = 1;cactus_sprite[1][10][66] = 1;cactus_sprite[1][10][67] = 1;cactus_sprite[1][10][68] = 1;cactus_sprite[1][10][69] = 1;cactus_sprite[1][11][34] = 1;cactus_sprite[1][11][35] = 1;cactus_sprite[1][11][36] = 1;cactus_sprite[1][11][37] = 1;cactus_sprite[1][11][38] = 1;cactus_sprite[1][11][39] = 1;cactus_sprite[1][11][40] = 1;cactus_sprite[1][11][41] = 1;cactus_sprite[1][11][42] = 1;cactus_sprite[1][11][43] = 1;cactus_sprite[1][11][44] = 1;cactus_sprite[1][11][45] = 1;cactus_sprite[1][11][46] = 1;cactus_sprite[1][11][47] = 1;cactus_sprite[1][11][48] = 1;cactus_sprite[1][11][49] = 1;cactus_sprite[1][11][50] = 1;cactus_sprite[1][11][51] = 1;cactus_sprite[1][11][52] = 1;cactus_sprite[1][11][53] = 1;cactus_sprite[1][11][54] = 1;cactus_sprite[1][11][55] = 1;cactus_sprite[1][11][56] = 1;cactus_sprite[1][11][57] = 1;cactus_sprite[1][11][58] = 1;cactus_sprite[1][11][59] = 1;cactus_sprite[1][11][60] = 1;cactus_sprite[1][11][61] = 1;cactus_sprite[1][11][62] = 1;cactus_sprite[1][11][63] = 1;cactus_sprite[1][11][64] = 1;cactus_sprite[1][11][65] = 1;cactus_sprite[1][11][66] = 1;cactus_sprite[1][11][67] = 1;cactus_sprite[1][11][68] = 1;cactus_sprite[1][11][69] = 1;cactus_sprite[1][12][60] = 1;cactus_sprite[1][12][61] = 1;cactus_sprite[1][12][62] = 1;cactus_sprite[1][12][63] = 1;cactus_sprite[1][12][64] = 1;cactus_sprite[1][12][65] = 1;cactus_sprite[1][12][66] = 1;cactus_sprite[1][12][67] = 1;cactus_sprite[1][12][68] = 1;cactus_sprite[1][12][69] = 1;cactus_sprite[1][13][60] = 1;cactus_sprite[1][13][61] = 1;cactus_sprite[1][13][62] = 1;cactus_sprite[1][13][63] = 1;cactus_sprite[1][13][64] = 1;cactus_sprite[1][13][65] = 1;cactus_sprite[1][13][66] = 1;cactus_sprite[1][13][67] = 1;cactus_sprite[1][13][68] = 1;cactus_sprite[1][13][69] = 1;cactus_sprite[1][14][60] = 1;cactus_sprite[1][14][61] = 1;cactus_sprite[1][14][62] = 1;cactus_sprite[1][14][63] = 1;cactus_sprite[1][14][64] = 1;cactus_sprite[1][14][65] = 1;cactus_sprite[1][14][66] = 1;cactus_sprite[1][14][67] = 1;cactus_sprite[1][14][68] = 1;cactus_sprite[1][14][69] = 1;cactus_sprite[1][15][60] = 1;cactus_sprite[1][15][61] = 1;cactus_sprite[1][15][62] = 1;cactus_sprite[1][15][63] = 1;cactus_sprite[1][15][64] = 1;cactus_sprite[1][15][65] = 1;cactus_sprite[1][15][66] = 1;cactus_sprite[1][15][67] = 1;cactus_sprite[1][15][68] = 1;cactus_sprite[1][15][69] = 1;cactus_sprite[1][16][60] = 1;cactus_sprite[1][16][61] = 1;cactus_sprite[1][16][62] = 1;cactus_sprite[1][16][63] = 1;cactus_sprite[1][16][64] = 1;cactus_sprite[1][16][65] = 1;cactus_sprite[1][16][66] = 1;cactus_sprite[1][16][67] = 1;cactus_sprite[1][16][68] = 1;cactus_sprite[1][16][69] = 1;cactus_sprite[1][17][60] = 1;cactus_sprite[1][17][61] = 1;cactus_sprite[1][17][62] = 1;cactus_sprite[1][17][63] = 1;cactus_sprite[1][17][64] = 1;cactus_sprite[1][17][65] = 1;cactus_sprite[1][17][66] = 1;cactus_sprite[1][17][67] = 1;cactus_sprite[1][17][68] = 1;cactus_sprite[1][17][69] = 1;cactus_sprite[1][18][10] = 1;cactus_sprite[1][18][11] = 1;cactus_sprite[1][18][12] = 1;cactus_sprite[1][18][13] = 1;cactus_sprite[1][18][14] = 1;cactus_sprite[1][18][15] = 1;cactus_sprite[1][18][16] = 1;cactus_sprite[1][18][17] = 1;cactus_sprite[1][18][18] = 1;cactus_sprite[1][18][19] = 1;cactus_sprite[1][18][20] = 1;cactus_sprite[1][18][21] = 1;cactus_sprite[1][18][22] = 1;cactus_sprite[1][18][23] = 1;cactus_sprite[1][18][24] = 1;cactus_sprite[1][18][25] = 1;cactus_sprite[1][18][26] = 1;cactus_sprite[1][18][27] = 1;cactus_sprite[1][18][28] = 1;cactus_sprite[1][18][29] = 1;cactus_sprite[1][18][30] = 1;cactus_sprite[1][18][31] = 1;cactus_sprite[1][18][32] = 1;cactus_sprite[1][18][33] = 1;cactus_sprite[1][18][34] = 1;cactus_sprite[1][18][35] = 1;cactus_sprite[1][18][36] = 1;cactus_sprite[1][18][37] = 1;cactus_sprite[1][18][38] = 1;cactus_sprite[1][18][39] = 1;cactus_sprite[1][18][40] = 1;cactus_sprite[1][18][41] = 1;cactus_sprite[1][18][42] = 1;cactus_sprite[1][18][43] = 1;cactus_sprite[1][18][44] = 1;cactus_sprite[1][18][45] = 1;cactus_sprite[1][18][46] = 1;cactus_sprite[1][18][47] = 1;cactus_sprite[1][18][48] = 1;cactus_sprite[1][18][49] = 1;cactus_sprite[1][18][50] = 1;cactus_sprite[1][18][51] = 1;cactus_sprite[1][18][52] = 1;cactus_sprite[1][18][53] = 1;cactus_sprite[1][18][54] = 1;cactus_sprite[1][18][55] = 1;cactus_sprite[1][18][56] = 1;cactus_sprite[1][18][57] = 1;cactus_sprite[1][18][58] = 1;cactus_sprite[1][18][59] = 1;cactus_sprite[1][18][60] = 1;cactus_sprite[1][18][61] = 1;cactus_sprite[1][18][62] = 1;cactus_sprite[1][18][63] = 1;cactus_sprite[1][18][64] = 1;cactus_sprite[1][18][65] = 1;cactus_sprite[1][18][66] = 1;cactus_sprite[1][18][67] = 1;cactus_sprite[1][18][68] = 1;cactus_sprite[1][18][69] = 1;cactus_sprite[1][18][70] = 1;cactus_sprite[1][18][71] = 1;cactus_sprite[1][18][72] = 1;cactus_sprite[1][18][73] = 1;cactus_sprite[1][18][74] = 1;cactus_sprite[1][18][75] = 1;cactus_sprite[1][18][76] = 1;cactus_sprite[1][18][77] = 1;cactus_sprite[1][18][78] = 1;cactus_sprite[1][18][79] = 1;cactus_sprite[1][18][80] = 1;cactus_sprite[1][18][81] = 1;cactus_sprite[1][18][82] = 1;cactus_sprite[1][18][83] = 1;cactus_sprite[1][18][84] = 1;cactus_sprite[1][18][85] = 1;cactus_sprite[1][18][86] = 1;cactus_sprite[1][18][87] = 1;cactus_sprite[1][18][88] = 1;cactus_sprite[1][18][89] = 1;cactus_sprite[1][18][90] = 1;cactus_sprite[1][18][91] = 1;cactus_sprite[1][18][92] = 1;cactus_sprite[1][18][93] = 1;cactus_sprite[1][18][94] = 1;cactus_sprite[1][18][95] = 1;cactus_sprite[1][18][96] = 1;cactus_sprite[1][18][97] = 1;cactus_sprite[1][18][98] = 1;cactus_sprite[1][18][99] = 1;cactus_sprite[1][19][10] = 1;cactus_sprite[1][19][11] = 1;cactus_sprite[1][19][12] = 1;cactus_sprite[1][19][13] = 1;cactus_sprite[1][19][14] = 1;cactus_sprite[1][19][15] = 1;cactus_sprite[1][19][16] = 1;cactus_sprite[1][19][17] = 1;cactus_sprite[1][19][18] = 1;cactus_sprite[1][19][19] = 1;cactus_sprite[1][19][20] = 1;cactus_sprite[1][19][21] = 1;cactus_sprite[1][19][22] = 1;cactus_sprite[1][19][23] = 1;cactus_sprite[1][19][24] = 1;cactus_sprite[1][19][25] = 1;cactus_sprite[1][19][26] = 1;cactus_sprite[1][19][27] = 1;cactus_sprite[1][19][28] = 1;cactus_sprite[1][19][29] = 1;cactus_sprite[1][19][30] = 1;cactus_sprite[1][19][31] = 1;cactus_sprite[1][19][32] = 1;cactus_sprite[1][19][33] = 1;cactus_sprite[1][19][34] = 1;cactus_sprite[1][19][35] = 1;cactus_sprite[1][19][36] = 1;cactus_sprite[1][19][37] = 1;cactus_sprite[1][19][38] = 1;cactus_sprite[1][19][39] = 1;cactus_sprite[1][19][40] = 1;cactus_sprite[1][19][41] = 1;cactus_sprite[1][19][42] = 1;cactus_sprite[1][19][43] = 1;cactus_sprite[1][19][44] = 1;cactus_sprite[1][19][45] = 1;cactus_sprite[1][19][46] = 1;cactus_sprite[1][19][47] = 1;cactus_sprite[1][19][48] = 1;cactus_sprite[1][19][49] = 1;cactus_sprite[1][19][50] = 1;cactus_sprite[1][19][51] = 1;cactus_sprite[1][19][52] = 1;cactus_sprite[1][19][53] = 1;cactus_sprite[1][19][54] = 1;cactus_sprite[1][19][55] = 1;cactus_sprite[1][19][56] = 1;cactus_sprite[1][19][57] = 1;cactus_sprite[1][19][58] = 1;cactus_sprite[1][19][59] = 1;cactus_sprite[1][19][60] = 1;cactus_sprite[1][19][61] = 1;cactus_sprite[1][19][62] = 1;cactus_sprite[1][19][63] = 1;cactus_sprite[1][19][64] = 1;cactus_sprite[1][19][65] = 1;cactus_sprite[1][19][66] = 1;cactus_sprite[1][19][67] = 1;cactus_sprite[1][19][68] = 1;cactus_sprite[1][19][69] = 1;cactus_sprite[1][19][70] = 1;cactus_sprite[1][19][71] = 1;cactus_sprite[1][19][72] = 1;cactus_sprite[1][19][73] = 1;cactus_sprite[1][19][74] = 1;cactus_sprite[1][19][75] = 1;cactus_sprite[1][19][76] = 1;cactus_sprite[1][19][77] = 1;cactus_sprite[1][19][78] = 1;cactus_sprite[1][19][79] = 1;cactus_sprite[1][19][80] = 1;cactus_sprite[1][19][81] = 1;cactus_sprite[1][19][82] = 1;cactus_sprite[1][19][83] = 1;cactus_sprite[1][19][84] = 1;cactus_sprite[1][19][85] = 1;cactus_sprite[1][19][86] = 1;cactus_sprite[1][19][87] = 1;cactus_sprite[1][19][88] = 1;cactus_sprite[1][19][89] = 1;cactus_sprite[1][19][90] = 1;cactus_sprite[1][19][91] = 1;cactus_sprite[1][19][92] = 1;cactus_sprite[1][19][93] = 1;cactus_sprite[1][19][94] = 1;cactus_sprite[1][19][95] = 1;cactus_sprite[1][19][96] = 1;cactus_sprite[1][19][97] = 1;cactus_sprite[1][19][98] = 1;cactus_sprite[1][19][99] = 1;cactus_sprite[1][20][8] = 1;cactus_sprite[1][20][9] = 1;cactus_sprite[1][20][10] = 1;cactus_sprite[1][20][11] = 1;cactus_sprite[1][20][12] = 1;cactus_sprite[1][20][13] = 1;cactus_sprite[1][20][14] = 1;cactus_sprite[1][20][15] = 1;cactus_sprite[1][20][16] = 1;cactus_sprite[1][20][17] = 1;cactus_sprite[1][20][18] = 1;cactus_sprite[1][20][19] = 1;cactus_sprite[1][20][20] = 1;cactus_sprite[1][20][21] = 1;cactus_sprite[1][20][22] = 1;cactus_sprite[1][20][23] = 1;cactus_sprite[1][20][24] = 1;cactus_sprite[1][20][25] = 1;cactus_sprite[1][20][26] = 1;cactus_sprite[1][20][27] = 1;cactus_sprite[1][20][28] = 1;cactus_sprite[1][20][29] = 1;cactus_sprite[1][20][30] = 1;cactus_sprite[1][20][31] = 1;cactus_sprite[1][20][32] = 1;cactus_sprite[1][20][33] = 1;cactus_sprite[1][20][34] = 1;cactus_sprite[1][20][35] = 1;cactus_sprite[1][20][36] = 1;cactus_sprite[1][20][37] = 1;cactus_sprite[1][20][38] = 1;cactus_sprite[1][20][39] = 1;cactus_sprite[1][20][40] = 1;cactus_sprite[1][20][41] = 1;cactus_sprite[1][20][42] = 1;cactus_sprite[1][20][43] = 1;cactus_sprite[1][20][44] = 1;cactus_sprite[1][20][45] = 1;cactus_sprite[1][20][46] = 1;cactus_sprite[1][20][47] = 1;cactus_sprite[1][20][48] = 1;cactus_sprite[1][20][49] = 1;cactus_sprite[1][20][50] = 1;cactus_sprite[1][20][51] = 1;cactus_sprite[1][20][52] = 1;cactus_sprite[1][20][53] = 1;cactus_sprite[1][20][54] = 1;cactus_sprite[1][20][55] = 1;cactus_sprite[1][20][56] = 1;cactus_sprite[1][20][57] = 1;cactus_sprite[1][20][58] = 1;cactus_sprite[1][20][59] = 1;cactus_sprite[1][20][60] = 1;cactus_sprite[1][20][61] = 1;cactus_sprite[1][20][62] = 1;cactus_sprite[1][20][63] = 1;cactus_sprite[1][20][64] = 1;cactus_sprite[1][20][65] = 1;cactus_sprite[1][20][66] = 1;cactus_sprite[1][20][67] = 1;cactus_sprite[1][20][68] = 1;cactus_sprite[1][20][69] = 1;cactus_sprite[1][20][70] = 1;cactus_sprite[1][20][71] = 1;cactus_sprite[1][20][72] = 1;cactus_sprite[1][20][73] = 1;cactus_sprite[1][20][74] = 1;cactus_sprite[1][20][75] = 1;cactus_sprite[1][20][76] = 1;cactus_sprite[1][20][77] = 1;cactus_sprite[1][20][78] = 1;cactus_sprite[1][20][79] = 1;cactus_sprite[1][20][80] = 1;cactus_sprite[1][20][81] = 1;cactus_sprite[1][20][82] = 1;cactus_sprite[1][20][83] = 1;cactus_sprite[1][20][84] = 1;cactus_sprite[1][20][85] = 1;cactus_sprite[1][20][86] = 1;cactus_sprite[1][20][87] = 1;cactus_sprite[1][20][88] = 1;cactus_sprite[1][20][89] = 1;cactus_sprite[1][20][90] = 1;cactus_sprite[1][20][91] = 1;cactus_sprite[1][20][92] = 1;cactus_sprite[1][20][93] = 1;cactus_sprite[1][20][94] = 1;cactus_sprite[1][20][95] = 1;cactus_sprite[1][20][96] = 1;cactus_sprite[1][20][97] = 1;cactus_sprite[1][20][98] = 1;cactus_sprite[1][20][99] = 1;cactus_sprite[1][21][8] = 1;cactus_sprite[1][21][9] = 1;cactus_sprite[1][21][10] = 1;cactus_sprite[1][21][11] = 1;cactus_sprite[1][21][12] = 1;cactus_sprite[1][21][13] = 1;cactus_sprite[1][21][14] = 1;cactus_sprite[1][21][15] = 1;cactus_sprite[1][21][16] = 1;cactus_sprite[1][21][17] = 1;cactus_sprite[1][21][18] = 1;cactus_sprite[1][21][19] = 1;cactus_sprite[1][21][20] = 1;cactus_sprite[1][21][21] = 1;cactus_sprite[1][21][22] = 1;cactus_sprite[1][21][23] = 1;cactus_sprite[1][21][24] = 1;cactus_sprite[1][21][25] = 1;cactus_sprite[1][21][26] = 1;cactus_sprite[1][21][27] = 1;cactus_sprite[1][21][28] = 1;cactus_sprite[1][21][29] = 1;cactus_sprite[1][21][30] = 1;cactus_sprite[1][21][31] = 1;cactus_sprite[1][21][32] = 1;cactus_sprite[1][21][33] = 1;cactus_sprite[1][21][34] = 1;cactus_sprite[1][21][35] = 1;cactus_sprite[1][21][36] = 1;cactus_sprite[1][21][37] = 1;cactus_sprite[1][21][38] = 1;cactus_sprite[1][21][39] = 1;cactus_sprite[1][21][40] = 1;cactus_sprite[1][21][41] = 1;cactus_sprite[1][21][42] = 1;cactus_sprite[1][21][43] = 1;cactus_sprite[1][21][44] = 1;cactus_sprite[1][21][45] = 1;cactus_sprite[1][21][46] = 1;cactus_sprite[1][21][47] = 1;cactus_sprite[1][21][48] = 1;cactus_sprite[1][21][49] = 1;cactus_sprite[1][21][50] = 1;cactus_sprite[1][21][51] = 1;cactus_sprite[1][21][52] = 1;cactus_sprite[1][21][53] = 1;cactus_sprite[1][21][54] = 1;cactus_sprite[1][21][55] = 1;cactus_sprite[1][21][56] = 1;cactus_sprite[1][21][57] = 1;cactus_sprite[1][21][58] = 1;cactus_sprite[1][21][59] = 1;cactus_sprite[1][21][60] = 1;cactus_sprite[1][21][61] = 1;cactus_sprite[1][21][62] = 1;cactus_sprite[1][21][63] = 1;cactus_sprite[1][21][64] = 1;cactus_sprite[1][21][65] = 1;cactus_sprite[1][21][66] = 1;cactus_sprite[1][21][67] = 1;cactus_sprite[1][21][68] = 1;cactus_sprite[1][21][69] = 1;cactus_sprite[1][21][70] = 1;cactus_sprite[1][21][71] = 1;cactus_sprite[1][21][72] = 1;cactus_sprite[1][21][73] = 1;cactus_sprite[1][21][74] = 1;cactus_sprite[1][21][75] = 1;cactus_sprite[1][21][76] = 1;cactus_sprite[1][21][77] = 1;cactus_sprite[1][21][78] = 1;cactus_sprite[1][21][79] = 1;cactus_sprite[1][21][80] = 1;cactus_sprite[1][21][81] = 1;cactus_sprite[1][21][82] = 1;cactus_sprite[1][21][83] = 1;cactus_sprite[1][21][84] = 1;cactus_sprite[1][21][85] = 1;cactus_sprite[1][21][86] = 1;cactus_sprite[1][21][87] = 1;cactus_sprite[1][21][88] = 1;cactus_sprite[1][21][89] = 1;cactus_sprite[1][21][90] = 1;cactus_sprite[1][21][91] = 1;cactus_sprite[1][21][92] = 1;cactus_sprite[1][21][93] = 1;cactus_sprite[1][21][94] = 1;cactus_sprite[1][21][95] = 1;cactus_sprite[1][21][96] = 1;cactus_sprite[1][21][97] = 1;cactus_sprite[1][21][98] = 1;cactus_sprite[1][21][99] = 1;cactus_sprite[1][22][8] = 1;cactus_sprite[1][22][9] = 1;cactus_sprite[1][22][10] = 1;cactus_sprite[1][22][11] = 1;cactus_sprite[1][22][12] = 1;cactus_sprite[1][22][13] = 1;cactus_sprite[1][22][14] = 1;cactus_sprite[1][22][15] = 1;cactus_sprite[1][22][16] = 1;cactus_sprite[1][22][17] = 1;cactus_sprite[1][22][18] = 1;cactus_sprite[1][22][19] = 1;cactus_sprite[1][22][20] = 1;cactus_sprite[1][22][21] = 1;cactus_sprite[1][22][22] = 1;cactus_sprite[1][22][23] = 1;cactus_sprite[1][22][24] = 1;cactus_sprite[1][22][25] = 1;cactus_sprite[1][22][26] = 1;cactus_sprite[1][22][27] = 1;cactus_sprite[1][22][28] = 1;cactus_sprite[1][22][29] = 1;cactus_sprite[1][22][30] = 1;cactus_sprite[1][22][31] = 1;cactus_sprite[1][22][32] = 1;cactus_sprite[1][22][33] = 1;cactus_sprite[1][22][34] = 1;cactus_sprite[1][22][35] = 1;cactus_sprite[1][22][36] = 1;cactus_sprite[1][22][37] = 1;cactus_sprite[1][22][38] = 1;cactus_sprite[1][22][39] = 1;cactus_sprite[1][22][40] = 1;cactus_sprite[1][22][41] = 1;cactus_sprite[1][22][42] = 1;cactus_sprite[1][22][43] = 1;cactus_sprite[1][22][44] = 1;cactus_sprite[1][22][45] = 1;cactus_sprite[1][22][46] = 1;cactus_sprite[1][22][47] = 1;cactus_sprite[1][22][48] = 1;cactus_sprite[1][22][49] = 1;cactus_sprite[1][22][50] = 1;cactus_sprite[1][22][51] = 1;cactus_sprite[1][22][52] = 1;cactus_sprite[1][22][53] = 1;cactus_sprite[1][22][54] = 1;cactus_sprite[1][22][55] = 1;cactus_sprite[1][22][56] = 1;cactus_sprite[1][22][57] = 1;cactus_sprite[1][22][58] = 1;cactus_sprite[1][22][59] = 1;cactus_sprite[1][22][60] = 1;cactus_sprite[1][22][61] = 1;cactus_sprite[1][22][62] = 1;cactus_sprite[1][22][63] = 1;cactus_sprite[1][22][64] = 1;cactus_sprite[1][22][65] = 1;cactus_sprite[1][22][66] = 1;cactus_sprite[1][22][67] = 1;cactus_sprite[1][22][68] = 1;cactus_sprite[1][22][69] = 1;cactus_sprite[1][22][70] = 1;cactus_sprite[1][22][71] = 1;cactus_sprite[1][22][72] = 1;cactus_sprite[1][22][73] = 1;cactus_sprite[1][22][74] = 1;cactus_sprite[1][22][75] = 1;cactus_sprite[1][22][76] = 1;cactus_sprite[1][22][77] = 1;cactus_sprite[1][22][78] = 1;cactus_sprite[1][22][79] = 1;cactus_sprite[1][22][80] = 1;cactus_sprite[1][22][81] = 1;cactus_sprite[1][22][82] = 1;cactus_sprite[1][22][83] = 1;cactus_sprite[1][22][84] = 1;cactus_sprite[1][22][85] = 1;cactus_sprite[1][22][86] = 1;cactus_sprite[1][22][87] = 1;cactus_sprite[1][22][88] = 1;cactus_sprite[1][22][89] = 1;cactus_sprite[1][22][90] = 1;cactus_sprite[1][22][91] = 1;cactus_sprite[1][22][92] = 1;cactus_sprite[1][22][93] = 1;cactus_sprite[1][22][94] = 1;cactus_sprite[1][22][95] = 1;cactus_sprite[1][22][96] = 1;cactus_sprite[1][22][97] = 1;cactus_sprite[1][22][98] = 1;cactus_sprite[1][22][99] = 1;cactus_sprite[1][23][8] = 1;cactus_sprite[1][23][9] = 1;cactus_sprite[1][23][10] = 1;cactus_sprite[1][23][11] = 1;cactus_sprite[1][23][12] = 1;cactus_sprite[1][23][13] = 1;cactus_sprite[1][23][14] = 1;cactus_sprite[1][23][15] = 1;cactus_sprite[1][23][16] = 1;cactus_sprite[1][23][17] = 1;cactus_sprite[1][23][18] = 1;cactus_sprite[1][23][19] = 1;cactus_sprite[1][23][20] = 1;cactus_sprite[1][23][21] = 1;cactus_sprite[1][23][22] = 1;cactus_sprite[1][23][23] = 1;cactus_sprite[1][23][24] = 1;cactus_sprite[1][23][25] = 1;cactus_sprite[1][23][26] = 1;cactus_sprite[1][23][27] = 1;cactus_sprite[1][23][28] = 1;cactus_sprite[1][23][29] = 1;cactus_sprite[1][23][30] = 1;cactus_sprite[1][23][31] = 1;cactus_sprite[1][23][32] = 1;cactus_sprite[1][23][33] = 1;cactus_sprite[1][23][34] = 1;cactus_sprite[1][23][35] = 1;cactus_sprite[1][23][36] = 1;cactus_sprite[1][23][37] = 1;cactus_sprite[1][23][38] = 1;cactus_sprite[1][23][39] = 1;cactus_sprite[1][23][40] = 1;cactus_sprite[1][23][41] = 1;cactus_sprite[1][23][42] = 1;cactus_sprite[1][23][43] = 1;cactus_sprite[1][23][44] = 1;cactus_sprite[1][23][45] = 1;cactus_sprite[1][23][46] = 1;cactus_sprite[1][23][47] = 1;cactus_sprite[1][23][48] = 1;cactus_sprite[1][23][49] = 1;cactus_sprite[1][23][50] = 1;cactus_sprite[1][23][51] = 1;cactus_sprite[1][23][52] = 1;cactus_sprite[1][23][53] = 1;cactus_sprite[1][23][54] = 1;cactus_sprite[1][23][55] = 1;cactus_sprite[1][23][56] = 1;cactus_sprite[1][23][57] = 1;cactus_sprite[1][23][58] = 1;cactus_sprite[1][23][59] = 1;cactus_sprite[1][23][60] = 1;cactus_sprite[1][23][61] = 1;cactus_sprite[1][23][62] = 1;cactus_sprite[1][23][63] = 1;cactus_sprite[1][23][64] = 1;cactus_sprite[1][23][65] = 1;cactus_sprite[1][23][66] = 1;cactus_sprite[1][23][67] = 1;cactus_sprite[1][23][68] = 1;cactus_sprite[1][23][69] = 1;cactus_sprite[1][23][70] = 1;cactus_sprite[1][23][71] = 1;cactus_sprite[1][23][72] = 1;cactus_sprite[1][23][73] = 1;cactus_sprite[1][23][74] = 1;cactus_sprite[1][23][75] = 1;cactus_sprite[1][23][76] = 1;cactus_sprite[1][23][77] = 1;cactus_sprite[1][23][78] = 1;cactus_sprite[1][23][79] = 1;cactus_sprite[1][23][80] = 1;cactus_sprite[1][23][81] = 1;cactus_sprite[1][23][82] = 1;cactus_sprite[1][23][83] = 1;cactus_sprite[1][23][84] = 1;cactus_sprite[1][23][85] = 1;cactus_sprite[1][23][86] = 1;cactus_sprite[1][23][87] = 1;cactus_sprite[1][23][88] = 1;cactus_sprite[1][23][89] = 1;cactus_sprite[1][23][90] = 1;cactus_sprite[1][23][91] = 1;cactus_sprite[1][23][92] = 1;cactus_sprite[1][23][93] = 1;cactus_sprite[1][23][94] = 1;cactus_sprite[1][23][95] = 1;cactus_sprite[1][23][96] = 1;cactus_sprite[1][23][97] = 1;cactus_sprite[1][23][98] = 1;cactus_sprite[1][23][99] = 1;cactus_sprite[1][24][8] = 1;cactus_sprite[1][24][9] = 1;cactus_sprite[1][24][10] = 1;cactus_sprite[1][24][11] = 1;cactus_sprite[1][24][12] = 1;cactus_sprite[1][24][13] = 1;cactus_sprite[1][24][14] = 1;cactus_sprite[1][24][15] = 1;cactus_sprite[1][24][16] = 1;cactus_sprite[1][24][17] = 1;cactus_sprite[1][24][18] = 1;cactus_sprite[1][24][19] = 1;cactus_sprite[1][24][20] = 1;cactus_sprite[1][24][21] = 1;cactus_sprite[1][24][22] = 1;cactus_sprite[1][24][23] = 1;cactus_sprite[1][24][24] = 1;cactus_sprite[1][24][25] = 1;cactus_sprite[1][24][26] = 1;cactus_sprite[1][24][27] = 1;cactus_sprite[1][24][28] = 1;cactus_sprite[1][24][29] = 1;cactus_sprite[1][24][30] = 1;cactus_sprite[1][24][31] = 1;cactus_sprite[1][24][32] = 1;cactus_sprite[1][24][33] = 1;cactus_sprite[1][24][34] = 1;cactus_sprite[1][24][35] = 1;cactus_sprite[1][24][36] = 1;cactus_sprite[1][24][37] = 1;cactus_sprite[1][24][38] = 1;cactus_sprite[1][24][39] = 1;cactus_sprite[1][24][40] = 1;cactus_sprite[1][24][41] = 1;cactus_sprite[1][24][42] = 1;cactus_sprite[1][24][43] = 1;cactus_sprite[1][24][44] = 1;cactus_sprite[1][24][45] = 1;cactus_sprite[1][24][46] = 1;cactus_sprite[1][24][47] = 1;cactus_sprite[1][24][48] = 1;cactus_sprite[1][24][49] = 1;cactus_sprite[1][24][50] = 1;cactus_sprite[1][24][51] = 1;cactus_sprite[1][24][52] = 1;cactus_sprite[1][24][53] = 1;cactus_sprite[1][24][54] = 1;cactus_sprite[1][24][55] = 1;cactus_sprite[1][24][56] = 1;cactus_sprite[1][24][57] = 1;cactus_sprite[1][24][58] = 1;cactus_sprite[1][24][59] = 1;cactus_sprite[1][24][60] = 1;cactus_sprite[1][24][61] = 1;cactus_sprite[1][24][62] = 1;cactus_sprite[1][24][63] = 1;cactus_sprite[1][24][64] = 1;cactus_sprite[1][24][65] = 1;cactus_sprite[1][24][66] = 1;cactus_sprite[1][24][67] = 1;cactus_sprite[1][24][68] = 1;cactus_sprite[1][24][69] = 1;cactus_sprite[1][24][70] = 1;cactus_sprite[1][24][71] = 1;cactus_sprite[1][24][72] = 1;cactus_sprite[1][24][73] = 1;cactus_sprite[1][24][74] = 1;cactus_sprite[1][24][75] = 1;cactus_sprite[1][24][76] = 1;cactus_sprite[1][24][77] = 1;cactus_sprite[1][24][78] = 1;cactus_sprite[1][24][79] = 1;cactus_sprite[1][24][80] = 1;cactus_sprite[1][24][81] = 1;cactus_sprite[1][24][82] = 1;cactus_sprite[1][24][83] = 1;cactus_sprite[1][24][84] = 1;cactus_sprite[1][24][85] = 1;cactus_sprite[1][24][86] = 1;cactus_sprite[1][24][87] = 1;cactus_sprite[1][24][88] = 1;cactus_sprite[1][24][89] = 1;cactus_sprite[1][24][90] = 1;cactus_sprite[1][24][91] = 1;cactus_sprite[1][24][92] = 1;cactus_sprite[1][24][93] = 1;cactus_sprite[1][24][94] = 1;cactus_sprite[1][24][95] = 1;cactus_sprite[1][24][96] = 1;cactus_sprite[1][24][97] = 1;cactus_sprite[1][24][98] = 1;cactus_sprite[1][24][99] = 1;cactus_sprite[1][25][8] = 1;cactus_sprite[1][25][9] = 1;cactus_sprite[1][25][10] = 1;cactus_sprite[1][25][11] = 1;cactus_sprite[1][25][12] = 1;cactus_sprite[1][25][13] = 1;cactus_sprite[1][25][14] = 1;cactus_sprite[1][25][15] = 1;cactus_sprite[1][25][16] = 1;cactus_sprite[1][25][17] = 1;cactus_sprite[1][25][18] = 1;cactus_sprite[1][25][19] = 1;cactus_sprite[1][25][20] = 1;cactus_sprite[1][25][21] = 1;cactus_sprite[1][25][22] = 1;cactus_sprite[1][25][23] = 1;cactus_sprite[1][25][24] = 1;cactus_sprite[1][25][25] = 1;cactus_sprite[1][25][26] = 1;cactus_sprite[1][25][27] = 1;cactus_sprite[1][25][28] = 1;cactus_sprite[1][25][29] = 1;cactus_sprite[1][25][30] = 1;cactus_sprite[1][25][31] = 1;cactus_sprite[1][25][32] = 1;cactus_sprite[1][25][33] = 1;cactus_sprite[1][25][34] = 1;cactus_sprite[1][25][35] = 1;cactus_sprite[1][25][36] = 1;cactus_sprite[1][25][37] = 1;cactus_sprite[1][25][38] = 1;cactus_sprite[1][25][39] = 1;cactus_sprite[1][25][40] = 1;cactus_sprite[1][25][41] = 1;cactus_sprite[1][25][42] = 1;cactus_sprite[1][25][43] = 1;cactus_sprite[1][25][44] = 1;cactus_sprite[1][25][45] = 1;cactus_sprite[1][25][46] = 1;cactus_sprite[1][25][47] = 1;cactus_sprite[1][25][48] = 1;cactus_sprite[1][25][49] = 1;cactus_sprite[1][25][50] = 1;cactus_sprite[1][25][51] = 1;cactus_sprite[1][25][52] = 1;cactus_sprite[1][25][53] = 1;cactus_sprite[1][25][54] = 1;cactus_sprite[1][25][55] = 1;cactus_sprite[1][25][56] = 1;cactus_sprite[1][25][57] = 1;cactus_sprite[1][25][58] = 1;cactus_sprite[1][25][59] = 1;cactus_sprite[1][25][60] = 1;cactus_sprite[1][25][61] = 1;cactus_sprite[1][25][62] = 1;cactus_sprite[1][25][63] = 1;cactus_sprite[1][25][64] = 1;cactus_sprite[1][25][65] = 1;cactus_sprite[1][25][66] = 1;cactus_sprite[1][25][67] = 1;cactus_sprite[1][25][68] = 1;cactus_sprite[1][25][69] = 1;cactus_sprite[1][25][70] = 1;cactus_sprite[1][25][71] = 1;cactus_sprite[1][25][72] = 1;cactus_sprite[1][25][73] = 1;cactus_sprite[1][25][74] = 1;cactus_sprite[1][25][75] = 1;cactus_sprite[1][25][76] = 1;cactus_sprite[1][25][77] = 1;cactus_sprite[1][25][78] = 1;cactus_sprite[1][25][79] = 1;cactus_sprite[1][25][80] = 1;cactus_sprite[1][25][81] = 1;cactus_sprite[1][25][82] = 1;cactus_sprite[1][25][83] = 1;cactus_sprite[1][25][84] = 1;cactus_sprite[1][25][85] = 1;cactus_sprite[1][25][86] = 1;cactus_sprite[1][25][87] = 1;cactus_sprite[1][25][88] = 1;cactus_sprite[1][25][89] = 1;cactus_sprite[1][25][90] = 1;cactus_sprite[1][25][91] = 1;cactus_sprite[1][25][92] = 1;cactus_sprite[1][25][93] = 1;cactus_sprite[1][25][94] = 1;cactus_sprite[1][25][95] = 1;cactus_sprite[1][25][96] = 1;cactus_sprite[1][25][97] = 1;cactus_sprite[1][25][98] = 1;cactus_sprite[1][25][99] = 1;cactus_sprite[1][26][8] = 1;cactus_sprite[1][26][9] = 1;cactus_sprite[1][26][10] = 1;cactus_sprite[1][26][11] = 1;cactus_sprite[1][26][12] = 1;cactus_sprite[1][26][13] = 1;cactus_sprite[1][26][14] = 1;cactus_sprite[1][26][15] = 1;cactus_sprite[1][26][16] = 1;cactus_sprite[1][26][17] = 1;cactus_sprite[1][26][18] = 1;cactus_sprite[1][26][19] = 1;cactus_sprite[1][26][20] = 1;cactus_sprite[1][26][21] = 1;cactus_sprite[1][26][22] = 1;cactus_sprite[1][26][23] = 1;cactus_sprite[1][26][24] = 1;cactus_sprite[1][26][25] = 1;cactus_sprite[1][26][26] = 1;cactus_sprite[1][26][27] = 1;cactus_sprite[1][26][28] = 1;cactus_sprite[1][26][29] = 1;cactus_sprite[1][26][30] = 1;cactus_sprite[1][26][31] = 1;cactus_sprite[1][26][32] = 1;cactus_sprite[1][26][33] = 1;cactus_sprite[1][26][34] = 1;cactus_sprite[1][26][35] = 1;cactus_sprite[1][26][36] = 1;cactus_sprite[1][26][37] = 1;cactus_sprite[1][26][38] = 1;cactus_sprite[1][26][39] = 1;cactus_sprite[1][26][40] = 1;cactus_sprite[1][26][41] = 1;cactus_sprite[1][26][42] = 1;cactus_sprite[1][26][43] = 1;cactus_sprite[1][26][44] = 1;cactus_sprite[1][26][45] = 1;cactus_sprite[1][26][46] = 1;cactus_sprite[1][26][47] = 1;cactus_sprite[1][26][48] = 1;cactus_sprite[1][26][49] = 1;cactus_sprite[1][26][50] = 1;cactus_sprite[1][26][51] = 1;cactus_sprite[1][26][52] = 1;cactus_sprite[1][26][53] = 1;cactus_sprite[1][26][54] = 1;cactus_sprite[1][26][55] = 1;cactus_sprite[1][26][56] = 1;cactus_sprite[1][26][57] = 1;cactus_sprite[1][26][58] = 1;cactus_sprite[1][26][59] = 1;cactus_sprite[1][26][60] = 1;cactus_sprite[1][26][61] = 1;cactus_sprite[1][26][62] = 1;cactus_sprite[1][26][63] = 1;cactus_sprite[1][26][64] = 1;cactus_sprite[1][26][65] = 1;cactus_sprite[1][26][66] = 1;cactus_sprite[1][26][67] = 1;cactus_sprite[1][26][68] = 1;cactus_sprite[1][26][69] = 1;cactus_sprite[1][26][70] = 1;cactus_sprite[1][26][71] = 1;cactus_sprite[1][26][72] = 1;cactus_sprite[1][26][73] = 1;cactus_sprite[1][26][74] = 1;cactus_sprite[1][26][75] = 1;cactus_sprite[1][26][76] = 1;cactus_sprite[1][26][77] = 1;cactus_sprite[1][26][78] = 1;cactus_sprite[1][26][79] = 1;cactus_sprite[1][26][80] = 1;cactus_sprite[1][26][81] = 1;cactus_sprite[1][26][82] = 1;cactus_sprite[1][26][83] = 1;cactus_sprite[1][26][84] = 1;cactus_sprite[1][26][85] = 1;cactus_sprite[1][26][86] = 1;cactus_sprite[1][26][87] = 1;cactus_sprite[1][26][88] = 1;cactus_sprite[1][26][89] = 1;cactus_sprite[1][26][90] = 1;cactus_sprite[1][26][91] = 1;cactus_sprite[1][26][92] = 1;cactus_sprite[1][26][93] = 1;cactus_sprite[1][26][94] = 1;cactus_sprite[1][26][95] = 1;cactus_sprite[1][26][96] = 1;cactus_sprite[1][26][97] = 1;cactus_sprite[1][26][98] = 1;cactus_sprite[1][26][99] = 1;cactus_sprite[1][27][8] = 1;cactus_sprite[1][27][9] = 1;cactus_sprite[1][27][10] = 1;cactus_sprite[1][27][11] = 1;cactus_sprite[1][27][12] = 1;cactus_sprite[1][27][13] = 1;cactus_sprite[1][27][14] = 1;cactus_sprite[1][27][15] = 1;cactus_sprite[1][27][16] = 1;cactus_sprite[1][27][17] = 1;cactus_sprite[1][27][18] = 1;cactus_sprite[1][27][19] = 1;cactus_sprite[1][27][20] = 1;cactus_sprite[1][27][21] = 1;cactus_sprite[1][27][22] = 1;cactus_sprite[1][27][23] = 1;cactus_sprite[1][27][24] = 1;cactus_sprite[1][27][25] = 1;cactus_sprite[1][27][26] = 1;cactus_sprite[1][27][27] = 1;cactus_sprite[1][27][28] = 1;cactus_sprite[1][27][29] = 1;cactus_sprite[1][27][30] = 1;cactus_sprite[1][27][31] = 1;cactus_sprite[1][27][32] = 1;cactus_sprite[1][27][33] = 1;cactus_sprite[1][27][34] = 1;cactus_sprite[1][27][35] = 1;cactus_sprite[1][27][36] = 1;cactus_sprite[1][27][37] = 1;cactus_sprite[1][27][38] = 1;cactus_sprite[1][27][39] = 1;cactus_sprite[1][27][40] = 1;cactus_sprite[1][27][41] = 1;cactus_sprite[1][27][42] = 1;cactus_sprite[1][27][43] = 1;cactus_sprite[1][27][44] = 1;cactus_sprite[1][27][45] = 1;cactus_sprite[1][27][46] = 1;cactus_sprite[1][27][47] = 1;cactus_sprite[1][27][48] = 1;cactus_sprite[1][27][49] = 1;cactus_sprite[1][27][50] = 1;cactus_sprite[1][27][51] = 1;cactus_sprite[1][27][52] = 1;cactus_sprite[1][27][53] = 1;cactus_sprite[1][27][54] = 1;cactus_sprite[1][27][55] = 1;cactus_sprite[1][27][56] = 1;cactus_sprite[1][27][57] = 1;cactus_sprite[1][27][58] = 1;cactus_sprite[1][27][59] = 1;cactus_sprite[1][27][60] = 1;cactus_sprite[1][27][61] = 1;cactus_sprite[1][27][62] = 1;cactus_sprite[1][27][63] = 1;cactus_sprite[1][27][64] = 1;cactus_sprite[1][27][65] = 1;cactus_sprite[1][27][66] = 1;cactus_sprite[1][27][67] = 1;cactus_sprite[1][27][68] = 1;cactus_sprite[1][27][69] = 1;cactus_sprite[1][27][70] = 1;cactus_sprite[1][27][71] = 1;cactus_sprite[1][27][72] = 1;cactus_sprite[1][27][73] = 1;cactus_sprite[1][27][74] = 1;cactus_sprite[1][27][75] = 1;cactus_sprite[1][27][76] = 1;cactus_sprite[1][27][77] = 1;cactus_sprite[1][27][78] = 1;cactus_sprite[1][27][79] = 1;cactus_sprite[1][27][80] = 1;cactus_sprite[1][27][81] = 1;cactus_sprite[1][27][82] = 1;cactus_sprite[1][27][83] = 1;cactus_sprite[1][27][84] = 1;cactus_sprite[1][27][85] = 1;cactus_sprite[1][27][86] = 1;cactus_sprite[1][27][87] = 1;cactus_sprite[1][27][88] = 1;cactus_sprite[1][27][89] = 1;cactus_sprite[1][27][90] = 1;cactus_sprite[1][27][91] = 1;cactus_sprite[1][27][92] = 1;cactus_sprite[1][27][93] = 1;cactus_sprite[1][27][94] = 1;cactus_sprite[1][27][95] = 1;cactus_sprite[1][27][96] = 1;cactus_sprite[1][27][97] = 1;cactus_sprite[1][27][98] = 1;cactus_sprite[1][27][99] = 1;cactus_sprite[1][28][8] = 1;cactus_sprite[1][28][9] = 1;cactus_sprite[1][28][10] = 1;cactus_sprite[1][28][11] = 1;cactus_sprite[1][28][12] = 1;cactus_sprite[1][28][13] = 1;cactus_sprite[1][28][14] = 1;cactus_sprite[1][28][15] = 1;cactus_sprite[1][28][16] = 1;cactus_sprite[1][28][17] = 1;cactus_sprite[1][28][18] = 1;cactus_sprite[1][28][19] = 1;cactus_sprite[1][28][20] = 1;cactus_sprite[1][28][21] = 1;cactus_sprite[1][28][22] = 1;cactus_sprite[1][28][23] = 1;cactus_sprite[1][28][24] = 1;cactus_sprite[1][28][25] = 1;cactus_sprite[1][28][26] = 1;cactus_sprite[1][28][27] = 1;cactus_sprite[1][28][28] = 1;cactus_sprite[1][28][29] = 1;cactus_sprite[1][28][30] = 1;cactus_sprite[1][28][31] = 1;cactus_sprite[1][28][32] = 1;cactus_sprite[1][28][33] = 1;cactus_sprite[1][28][34] = 1;cactus_sprite[1][28][35] = 1;cactus_sprite[1][28][36] = 1;cactus_sprite[1][28][37] = 1;cactus_sprite[1][28][38] = 1;cactus_sprite[1][28][39] = 1;cactus_sprite[1][28][40] = 1;cactus_sprite[1][28][41] = 1;cactus_sprite[1][28][42] = 1;cactus_sprite[1][28][43] = 1;cactus_sprite[1][28][44] = 1;cactus_sprite[1][28][45] = 1;cactus_sprite[1][28][46] = 1;cactus_sprite[1][28][47] = 1;cactus_sprite[1][28][48] = 1;cactus_sprite[1][28][49] = 1;cactus_sprite[1][28][50] = 1;cactus_sprite[1][28][51] = 1;cactus_sprite[1][28][52] = 1;cactus_sprite[1][28][53] = 1;cactus_sprite[1][28][54] = 1;cactus_sprite[1][28][55] = 1;cactus_sprite[1][28][56] = 1;cactus_sprite[1][28][57] = 1;cactus_sprite[1][28][58] = 1;cactus_sprite[1][28][59] = 1;cactus_sprite[1][28][60] = 1;cactus_sprite[1][28][61] = 1;cactus_sprite[1][28][62] = 1;cactus_sprite[1][28][63] = 1;cactus_sprite[1][28][64] = 1;cactus_sprite[1][28][65] = 1;cactus_sprite[1][28][66] = 1;cactus_sprite[1][28][67] = 1;cactus_sprite[1][28][68] = 1;cactus_sprite[1][28][69] = 1;cactus_sprite[1][28][70] = 1;cactus_sprite[1][28][71] = 1;cactus_sprite[1][28][72] = 1;cactus_sprite[1][28][73] = 1;cactus_sprite[1][28][74] = 1;cactus_sprite[1][28][75] = 1;cactus_sprite[1][28][76] = 1;cactus_sprite[1][28][77] = 1;cactus_sprite[1][28][78] = 1;cactus_sprite[1][28][79] = 1;cactus_sprite[1][28][80] = 1;cactus_sprite[1][28][81] = 1;cactus_sprite[1][28][82] = 1;cactus_sprite[1][28][83] = 1;cactus_sprite[1][28][84] = 1;cactus_sprite[1][28][85] = 1;cactus_sprite[1][28][86] = 1;cactus_sprite[1][28][87] = 1;cactus_sprite[1][28][88] = 1;cactus_sprite[1][28][89] = 1;cactus_sprite[1][28][90] = 1;cactus_sprite[1][28][91] = 1;cactus_sprite[1][28][92] = 1;cactus_sprite[1][28][93] = 1;cactus_sprite[1][28][94] = 1;cactus_sprite[1][28][95] = 1;cactus_sprite[1][28][96] = 1;cactus_sprite[1][28][97] = 1;cactus_sprite[1][28][98] = 1;cactus_sprite[1][28][99] = 1;cactus_sprite[1][29][8] = 1;cactus_sprite[1][29][9] = 1;cactus_sprite[1][29][10] = 1;cactus_sprite[1][29][11] = 1;cactus_sprite[1][29][12] = 1;cactus_sprite[1][29][13] = 1;cactus_sprite[1][29][14] = 1;cactus_sprite[1][29][15] = 1;cactus_sprite[1][29][16] = 1;cactus_sprite[1][29][17] = 1;cactus_sprite[1][29][18] = 1;cactus_sprite[1][29][19] = 1;cactus_sprite[1][29][20] = 1;cactus_sprite[1][29][21] = 1;cactus_sprite[1][29][22] = 1;cactus_sprite[1][29][23] = 1;cactus_sprite[1][29][24] = 1;cactus_sprite[1][29][25] = 1;cactus_sprite[1][29][26] = 1;cactus_sprite[1][29][27] = 1;cactus_sprite[1][29][28] = 1;cactus_sprite[1][29][29] = 1;cactus_sprite[1][29][30] = 1;cactus_sprite[1][29][31] = 1;cactus_sprite[1][29][32] = 1;cactus_sprite[1][29][33] = 1;cactus_sprite[1][29][34] = 1;cactus_sprite[1][29][35] = 1;cactus_sprite[1][29][36] = 1;cactus_sprite[1][29][37] = 1;cactus_sprite[1][29][38] = 1;cactus_sprite[1][29][39] = 1;cactus_sprite[1][29][40] = 1;cactus_sprite[1][29][41] = 1;cactus_sprite[1][29][42] = 1;cactus_sprite[1][29][43] = 1;cactus_sprite[1][29][44] = 1;cactus_sprite[1][29][45] = 1;cactus_sprite[1][29][46] = 1;cactus_sprite[1][29][47] = 1;cactus_sprite[1][29][48] = 1;cactus_sprite[1][29][49] = 1;cactus_sprite[1][29][50] = 1;cactus_sprite[1][29][51] = 1;cactus_sprite[1][29][52] = 1;cactus_sprite[1][29][53] = 1;cactus_sprite[1][29][54] = 1;cactus_sprite[1][29][55] = 1;cactus_sprite[1][29][56] = 1;cactus_sprite[1][29][57] = 1;cactus_sprite[1][29][58] = 1;cactus_sprite[1][29][59] = 1;cactus_sprite[1][29][60] = 1;cactus_sprite[1][29][61] = 1;cactus_sprite[1][29][62] = 1;cactus_sprite[1][29][63] = 1;cactus_sprite[1][29][64] = 1;cactus_sprite[1][29][65] = 1;cactus_sprite[1][29][66] = 1;cactus_sprite[1][29][67] = 1;cactus_sprite[1][29][68] = 1;cactus_sprite[1][29][69] = 1;cactus_sprite[1][29][70] = 1;cactus_sprite[1][29][71] = 1;cactus_sprite[1][29][72] = 1;cactus_sprite[1][29][73] = 1;cactus_sprite[1][29][74] = 1;cactus_sprite[1][29][75] = 1;cactus_sprite[1][29][76] = 1;cactus_sprite[1][29][77] = 1;cactus_sprite[1][29][78] = 1;cactus_sprite[1][29][79] = 1;cactus_sprite[1][29][80] = 1;cactus_sprite[1][29][81] = 1;cactus_sprite[1][29][82] = 1;cactus_sprite[1][29][83] = 1;cactus_sprite[1][29][84] = 1;cactus_sprite[1][29][85] = 1;cactus_sprite[1][29][86] = 1;cactus_sprite[1][29][87] = 1;cactus_sprite[1][29][88] = 1;cactus_sprite[1][29][89] = 1;cactus_sprite[1][29][90] = 1;cactus_sprite[1][29][91] = 1;cactus_sprite[1][29][92] = 1;cactus_sprite[1][29][93] = 1;cactus_sprite[1][29][94] = 1;cactus_sprite[1][29][95] = 1;cactus_sprite[1][29][96] = 1;cactus_sprite[1][29][97] = 1;cactus_sprite[1][29][98] = 1;cactus_sprite[1][29][99] = 1;cactus_sprite[1][30][10] = 1;cactus_sprite[1][30][11] = 1;cactus_sprite[1][30][12] = 1;cactus_sprite[1][30][13] = 1;cactus_sprite[1][30][14] = 1;cactus_sprite[1][30][15] = 1;cactus_sprite[1][30][16] = 1;cactus_sprite[1][30][17] = 1;cactus_sprite[1][30][18] = 1;cactus_sprite[1][30][19] = 1;cactus_sprite[1][30][20] = 1;cactus_sprite[1][30][21] = 1;cactus_sprite[1][30][22] = 1;cactus_sprite[1][30][23] = 1;cactus_sprite[1][30][24] = 1;cactus_sprite[1][30][25] = 1;cactus_sprite[1][30][26] = 1;cactus_sprite[1][30][27] = 1;cactus_sprite[1][30][28] = 1;cactus_sprite[1][30][29] = 1;cactus_sprite[1][30][30] = 1;cactus_sprite[1][30][31] = 1;cactus_sprite[1][30][32] = 1;cactus_sprite[1][30][33] = 1;cactus_sprite[1][30][34] = 1;cactus_sprite[1][30][35] = 1;cactus_sprite[1][30][36] = 1;cactus_sprite[1][30][37] = 1;cactus_sprite[1][30][38] = 1;cactus_sprite[1][30][39] = 1;cactus_sprite[1][30][40] = 1;cactus_sprite[1][30][41] = 1;cactus_sprite[1][30][42] = 1;cactus_sprite[1][30][43] = 1;cactus_sprite[1][30][44] = 1;cactus_sprite[1][30][45] = 1;cactus_sprite[1][30][46] = 1;cactus_sprite[1][30][47] = 1;cactus_sprite[1][30][48] = 1;cactus_sprite[1][30][49] = 1;cactus_sprite[1][30][50] = 1;cactus_sprite[1][30][51] = 1;cactus_sprite[1][30][52] = 1;cactus_sprite[1][30][53] = 1;cactus_sprite[1][30][54] = 1;cactus_sprite[1][30][55] = 1;cactus_sprite[1][30][56] = 1;cactus_sprite[1][30][57] = 1;cactus_sprite[1][30][58] = 1;cactus_sprite[1][30][59] = 1;cactus_sprite[1][30][60] = 1;cactus_sprite[1][30][61] = 1;cactus_sprite[1][30][62] = 1;cactus_sprite[1][30][63] = 1;cactus_sprite[1][30][64] = 1;cactus_sprite[1][30][65] = 1;cactus_sprite[1][30][66] = 1;cactus_sprite[1][30][67] = 1;cactus_sprite[1][30][68] = 1;cactus_sprite[1][30][69] = 1;cactus_sprite[1][30][70] = 1;cactus_sprite[1][30][71] = 1;cactus_sprite[1][30][72] = 1;cactus_sprite[1][30][73] = 1;cactus_sprite[1][30][74] = 1;cactus_sprite[1][30][75] = 1;cactus_sprite[1][30][76] = 1;cactus_sprite[1][30][77] = 1;cactus_sprite[1][30][78] = 1;cactus_sprite[1][30][79] = 1;cactus_sprite[1][30][80] = 1;cactus_sprite[1][30][81] = 1;cactus_sprite[1][30][82] = 1;cactus_sprite[1][30][83] = 1;cactus_sprite[1][30][84] = 1;cactus_sprite[1][30][85] = 1;cactus_sprite[1][30][86] = 1;cactus_sprite[1][30][87] = 1;cactus_sprite[1][30][88] = 1;cactus_sprite[1][30][89] = 1;cactus_sprite[1][30][90] = 1;cactus_sprite[1][30][91] = 1;cactus_sprite[1][30][92] = 1;cactus_sprite[1][30][93] = 1;cactus_sprite[1][30][94] = 1;cactus_sprite[1][30][95] = 1;cactus_sprite[1][30][96] = 1;cactus_sprite[1][30][97] = 1;cactus_sprite[1][30][98] = 1;cactus_sprite[1][30][99] = 1;cactus_sprite[1][31][10] = 1;cactus_sprite[1][31][11] = 1;cactus_sprite[1][31][12] = 1;cactus_sprite[1][31][13] = 1;cactus_sprite[1][31][14] = 1;cactus_sprite[1][31][15] = 1;cactus_sprite[1][31][16] = 1;cactus_sprite[1][31][17] = 1;cactus_sprite[1][31][18] = 1;cactus_sprite[1][31][19] = 1;cactus_sprite[1][31][20] = 1;cactus_sprite[1][31][21] = 1;cactus_sprite[1][31][22] = 1;cactus_sprite[1][31][23] = 1;cactus_sprite[1][31][24] = 1;cactus_sprite[1][31][25] = 1;cactus_sprite[1][31][26] = 1;cactus_sprite[1][31][27] = 1;cactus_sprite[1][31][28] = 1;cactus_sprite[1][31][29] = 1;cactus_sprite[1][31][30] = 1;cactus_sprite[1][31][31] = 1;cactus_sprite[1][31][32] = 1;cactus_sprite[1][31][33] = 1;cactus_sprite[1][31][34] = 1;cactus_sprite[1][31][35] = 1;cactus_sprite[1][31][36] = 1;cactus_sprite[1][31][37] = 1;cactus_sprite[1][31][38] = 1;cactus_sprite[1][31][39] = 1;cactus_sprite[1][31][40] = 1;cactus_sprite[1][31][41] = 1;cactus_sprite[1][31][42] = 1;cactus_sprite[1][31][43] = 1;cactus_sprite[1][31][44] = 1;cactus_sprite[1][31][45] = 1;cactus_sprite[1][31][46] = 1;cactus_sprite[1][31][47] = 1;cactus_sprite[1][31][48] = 1;cactus_sprite[1][31][49] = 1;cactus_sprite[1][31][50] = 1;cactus_sprite[1][31][51] = 1;cactus_sprite[1][31][52] = 1;cactus_sprite[1][31][53] = 1;cactus_sprite[1][31][54] = 1;cactus_sprite[1][31][55] = 1;cactus_sprite[1][31][56] = 1;cactus_sprite[1][31][57] = 1;cactus_sprite[1][31][58] = 1;cactus_sprite[1][31][59] = 1;cactus_sprite[1][31][60] = 1;cactus_sprite[1][31][61] = 1;cactus_sprite[1][31][62] = 1;cactus_sprite[1][31][63] = 1;cactus_sprite[1][31][64] = 1;cactus_sprite[1][31][65] = 1;cactus_sprite[1][31][66] = 1;cactus_sprite[1][31][67] = 1;cactus_sprite[1][31][68] = 1;cactus_sprite[1][31][69] = 1;cactus_sprite[1][31][70] = 1;cactus_sprite[1][31][71] = 1;cactus_sprite[1][31][72] = 1;cactus_sprite[1][31][73] = 1;cactus_sprite[1][31][74] = 1;cactus_sprite[1][31][75] = 1;cactus_sprite[1][31][76] = 1;cactus_sprite[1][31][77] = 1;cactus_sprite[1][31][78] = 1;cactus_sprite[1][31][79] = 1;cactus_sprite[1][31][80] = 1;cactus_sprite[1][31][81] = 1;cactus_sprite[1][31][82] = 1;cactus_sprite[1][31][83] = 1;cactus_sprite[1][31][84] = 1;cactus_sprite[1][31][85] = 1;cactus_sprite[1][31][86] = 1;cactus_sprite[1][31][87] = 1;cactus_sprite[1][31][88] = 1;cactus_sprite[1][31][89] = 1;cactus_sprite[1][31][90] = 1;cactus_sprite[1][31][91] = 1;cactus_sprite[1][31][92] = 1;cactus_sprite[1][31][93] = 1;cactus_sprite[1][31][94] = 1;cactus_sprite[1][31][95] = 1;cactus_sprite[1][31][96] = 1;cactus_sprite[1][31][97] = 1;cactus_sprite[1][31][98] = 1;cactus_sprite[1][31][99] = 1;cactus_sprite[1][32][60] = 1;cactus_sprite[1][32][61] = 1;cactus_sprite[1][32][62] = 1;cactus_sprite[1][32][63] = 1;cactus_sprite[1][32][64] = 1;cactus_sprite[1][32][65] = 1;cactus_sprite[1][32][66] = 1;cactus_sprite[1][32][67] = 1;cactus_sprite[1][33][60] = 1;cactus_sprite[1][33][61] = 1;cactus_sprite[1][33][62] = 1;cactus_sprite[1][33][63] = 1;cactus_sprite[1][33][64] = 1;cactus_sprite[1][33][65] = 1;cactus_sprite[1][33][66] = 1;cactus_sprite[1][33][67] = 1;cactus_sprite[1][34][60] = 1;cactus_sprite[1][34][61] = 1;cactus_sprite[1][34][62] = 1;cactus_sprite[1][34][63] = 1;cactus_sprite[1][34][64] = 1;cactus_sprite[1][34][65] = 1;cactus_sprite[1][34][66] = 1;cactus_sprite[1][34][67] = 1;cactus_sprite[1][35][60] = 1;cactus_sprite[1][35][61] = 1;cactus_sprite[1][35][62] = 1;cactus_sprite[1][35][63] = 1;cactus_sprite[1][35][64] = 1;cactus_sprite[1][35][65] = 1;cactus_sprite[1][35][66] = 1;cactus_sprite[1][35][67] = 1;cactus_sprite[1][36][60] = 1;cactus_sprite[1][36][61] = 1;cactus_sprite[1][36][62] = 1;cactus_sprite[1][36][63] = 1;cactus_sprite[1][36][64] = 1;cactus_sprite[1][36][65] = 1;cactus_sprite[1][36][66] = 1;cactus_sprite[1][36][67] = 1;cactus_sprite[1][37][60] = 1;cactus_sprite[1][37][61] = 1;cactus_sprite[1][37][62] = 1;cactus_sprite[1][37][63] = 1;cactus_sprite[1][37][64] = 1;cactus_sprite[1][37][65] = 1;cactus_sprite[1][37][66] = 1;cactus_sprite[1][37][67] = 1;cactus_sprite[1][38][30] = 1;cactus_sprite[1][38][31] = 1;cactus_sprite[1][38][32] = 1;cactus_sprite[1][38][33] = 1;cactus_sprite[1][38][34] = 1;cactus_sprite[1][38][35] = 1;cactus_sprite[1][38][36] = 1;cactus_sprite[1][38][37] = 1;cactus_sprite[1][38][38] = 1;cactus_sprite[1][38][39] = 1;cactus_sprite[1][38][40] = 1;cactus_sprite[1][38][41] = 1;cactus_sprite[1][38][42] = 1;cactus_sprite[1][38][43] = 1;cactus_sprite[1][38][44] = 1;cactus_sprite[1][38][45] = 1;cactus_sprite[1][38][46] = 1;cactus_sprite[1][38][47] = 1;cactus_sprite[1][38][48] = 1;cactus_sprite[1][38][49] = 1;cactus_sprite[1][38][50] = 1;cactus_sprite[1][38][51] = 1;cactus_sprite[1][38][52] = 1;cactus_sprite[1][38][53] = 1;cactus_sprite[1][38][54] = 1;cactus_sprite[1][38][55] = 1;cactus_sprite[1][38][56] = 1;cactus_sprite[1][38][57] = 1;cactus_sprite[1][38][58] = 1;cactus_sprite[1][38][59] = 1;cactus_sprite[1][38][60] = 1;cactus_sprite[1][38][61] = 1;cactus_sprite[1][38][62] = 1;cactus_sprite[1][38][63] = 1;cactus_sprite[1][38][64] = 1;cactus_sprite[1][38][65] = 1;cactus_sprite[1][38][66] = 1;cactus_sprite[1][38][67] = 1;cactus_sprite[1][39][30] = 1;cactus_sprite[1][39][31] = 1;cactus_sprite[1][39][32] = 1;cactus_sprite[1][39][33] = 1;cactus_sprite[1][39][34] = 1;cactus_sprite[1][39][35] = 1;cactus_sprite[1][39][36] = 1;cactus_sprite[1][39][37] = 1;cactus_sprite[1][39][38] = 1;cactus_sprite[1][39][39] = 1;cactus_sprite[1][39][40] = 1;cactus_sprite[1][39][41] = 1;cactus_sprite[1][39][42] = 1;cactus_sprite[1][39][43] = 1;cactus_sprite[1][39][44] = 1;cactus_sprite[1][39][45] = 1;cactus_sprite[1][39][46] = 1;cactus_sprite[1][39][47] = 1;cactus_sprite[1][39][48] = 1;cactus_sprite[1][39][49] = 1;cactus_sprite[1][39][50] = 1;cactus_sprite[1][39][51] = 1;cactus_sprite[1][39][52] = 1;cactus_sprite[1][39][53] = 1;cactus_sprite[1][39][54] = 1;cactus_sprite[1][39][55] = 1;cactus_sprite[1][39][56] = 1;cactus_sprite[1][39][57] = 1;cactus_sprite[1][39][58] = 1;cactus_sprite[1][39][59] = 1;cactus_sprite[1][39][60] = 1;cactus_sprite[1][39][61] = 1;cactus_sprite[1][39][62] = 1;cactus_sprite[1][39][63] = 1;cactus_sprite[1][39][64] = 1;cactus_sprite[1][39][65] = 1;cactus_sprite[1][39][66] = 1;cactus_sprite[1][39][67] = 1;cactus_sprite[1][40][28] = 1;cactus_sprite[1][40][29] = 1;cactus_sprite[1][40][30] = 1;cactus_sprite[1][40][31] = 1;cactus_sprite[1][40][32] = 1;cactus_sprite[1][40][33] = 1;cactus_sprite[1][40][34] = 1;cactus_sprite[1][40][35] = 1;cactus_sprite[1][40][36] = 1;cactus_sprite[1][40][37] = 1;cactus_sprite[1][40][38] = 1;cactus_sprite[1][40][39] = 1;cactus_sprite[1][40][40] = 1;cactus_sprite[1][40][41] = 1;cactus_sprite[1][40][42] = 1;cactus_sprite[1][40][43] = 1;cactus_sprite[1][40][44] = 1;cactus_sprite[1][40][45] = 1;cactus_sprite[1][40][46] = 1;cactus_sprite[1][40][47] = 1;cactus_sprite[1][40][48] = 1;cactus_sprite[1][40][49] = 1;cactus_sprite[1][40][50] = 1;cactus_sprite[1][40][51] = 1;cactus_sprite[1][40][52] = 1;cactus_sprite[1][40][53] = 1;cactus_sprite[1][40][54] = 1;cactus_sprite[1][40][55] = 1;cactus_sprite[1][40][56] = 1;cactus_sprite[1][40][57] = 1;cactus_sprite[1][40][58] = 1;cactus_sprite[1][40][59] = 1;cactus_sprite[1][40][60] = 1;cactus_sprite[1][40][61] = 1;cactus_sprite[1][40][62] = 1;cactus_sprite[1][40][63] = 1;cactus_sprite[1][40][64] = 1;cactus_sprite[1][40][65] = 1;cactus_sprite[1][41][28] = 1;cactus_sprite[1][41][29] = 1;cactus_sprite[1][41][30] = 1;cactus_sprite[1][41][31] = 1;cactus_sprite[1][41][32] = 1;cactus_sprite[1][41][33] = 1;cactus_sprite[1][41][34] = 1;cactus_sprite[1][41][35] = 1;cactus_sprite[1][41][36] = 1;cactus_sprite[1][41][37] = 1;cactus_sprite[1][41][38] = 1;cactus_sprite[1][41][39] = 1;cactus_sprite[1][41][40] = 1;cactus_sprite[1][41][41] = 1;cactus_sprite[1][41][42] = 1;cactus_sprite[1][41][43] = 1;cactus_sprite[1][41][44] = 1;cactus_sprite[1][41][45] = 1;cactus_sprite[1][41][46] = 1;cactus_sprite[1][41][47] = 1;cactus_sprite[1][41][48] = 1;cactus_sprite[1][41][49] = 1;cactus_sprite[1][41][50] = 1;cactus_sprite[1][41][51] = 1;cactus_sprite[1][41][52] = 1;cactus_sprite[1][41][53] = 1;cactus_sprite[1][41][54] = 1;cactus_sprite[1][41][55] = 1;cactus_sprite[1][41][56] = 1;cactus_sprite[1][41][57] = 1;cactus_sprite[1][41][58] = 1;cactus_sprite[1][41][59] = 1;cactus_sprite[1][41][60] = 1;cactus_sprite[1][41][61] = 1;cactus_sprite[1][41][62] = 1;cactus_sprite[1][41][63] = 1;cactus_sprite[1][41][64] = 1;cactus_sprite[1][41][65] = 1;cactus_sprite[1][42][28] = 1;cactus_sprite[1][42][29] = 1;cactus_sprite[1][42][30] = 1;cactus_sprite[1][42][31] = 1;cactus_sprite[1][42][32] = 1;cactus_sprite[1][42][33] = 1;cactus_sprite[1][42][34] = 1;cactus_sprite[1][42][35] = 1;cactus_sprite[1][42][36] = 1;cactus_sprite[1][42][37] = 1;cactus_sprite[1][42][38] = 1;cactus_sprite[1][42][39] = 1;cactus_sprite[1][42][40] = 1;cactus_sprite[1][42][41] = 1;cactus_sprite[1][42][42] = 1;cactus_sprite[1][42][43] = 1;cactus_sprite[1][42][44] = 1;cactus_sprite[1][42][45] = 1;cactus_sprite[1][42][46] = 1;cactus_sprite[1][42][47] = 1;cactus_sprite[1][42][48] = 1;cactus_sprite[1][42][49] = 1;cactus_sprite[1][42][50] = 1;cactus_sprite[1][42][51] = 1;cactus_sprite[1][42][52] = 1;cactus_sprite[1][42][53] = 1;cactus_sprite[1][42][54] = 1;cactus_sprite[1][42][55] = 1;cactus_sprite[1][42][56] = 1;cactus_sprite[1][42][57] = 1;cactus_sprite[1][42][58] = 1;cactus_sprite[1][42][59] = 1;cactus_sprite[1][42][60] = 1;cactus_sprite[1][42][61] = 1;cactus_sprite[1][42][62] = 1;cactus_sprite[1][42][63] = 1;cactus_sprite[1][43][28] = 1;cactus_sprite[1][43][29] = 1;cactus_sprite[1][43][30] = 1;cactus_sprite[1][43][31] = 1;cactus_sprite[1][43][32] = 1;cactus_sprite[1][43][33] = 1;cactus_sprite[1][43][34] = 1;cactus_sprite[1][43][35] = 1;cactus_sprite[1][43][36] = 1;cactus_sprite[1][43][37] = 1;cactus_sprite[1][43][38] = 1;cactus_sprite[1][43][39] = 1;cactus_sprite[1][43][40] = 1;cactus_sprite[1][43][41] = 1;cactus_sprite[1][43][42] = 1;cactus_sprite[1][43][43] = 1;cactus_sprite[1][43][44] = 1;cactus_sprite[1][43][45] = 1;cactus_sprite[1][43][46] = 1;cactus_sprite[1][43][47] = 1;cactus_sprite[1][43][48] = 1;cactus_sprite[1][43][49] = 1;cactus_sprite[1][43][50] = 1;cactus_sprite[1][43][51] = 1;cactus_sprite[1][43][52] = 1;cactus_sprite[1][43][53] = 1;cactus_sprite[1][43][54] = 1;cactus_sprite[1][43][55] = 1;cactus_sprite[1][43][56] = 1;cactus_sprite[1][43][57] = 1;cactus_sprite[1][43][58] = 1;cactus_sprite[1][43][59] = 1;cactus_sprite[1][43][60] = 1;cactus_sprite[1][43][61] = 1;cactus_sprite[1][43][62] = 1;cactus_sprite[1][43][63] = 1;cactus_sprite[1][44][28] = 1;cactus_sprite[1][44][29] = 1;cactus_sprite[1][44][30] = 1;cactus_sprite[1][44][31] = 1;cactus_sprite[1][44][32] = 1;cactus_sprite[1][44][33] = 1;cactus_sprite[1][44][34] = 1;cactus_sprite[1][44][35] = 1;cactus_sprite[1][44][36] = 1;cactus_sprite[1][44][37] = 1;cactus_sprite[1][44][38] = 1;cactus_sprite[1][44][39] = 1;cactus_sprite[1][44][40] = 1;cactus_sprite[1][44][41] = 1;cactus_sprite[1][44][42] = 1;cactus_sprite[1][44][43] = 1;cactus_sprite[1][44][44] = 1;cactus_sprite[1][44][45] = 1;cactus_sprite[1][44][46] = 1;cactus_sprite[1][44][47] = 1;cactus_sprite[1][44][48] = 1;cactus_sprite[1][44][49] = 1;cactus_sprite[1][44][50] = 1;cactus_sprite[1][44][51] = 1;cactus_sprite[1][44][52] = 1;cactus_sprite[1][44][53] = 1;cactus_sprite[1][44][54] = 1;cactus_sprite[1][44][55] = 1;cactus_sprite[1][44][56] = 1;cactus_sprite[1][44][57] = 1;cactus_sprite[1][44][58] = 1;cactus_sprite[1][44][59] = 1;cactus_sprite[1][44][60] = 1;cactus_sprite[1][44][61] = 1;cactus_sprite[1][45][28] = 1;cactus_sprite[1][45][29] = 1;cactus_sprite[1][45][30] = 1;cactus_sprite[1][45][31] = 1;cactus_sprite[1][45][32] = 1;cactus_sprite[1][45][33] = 1;cactus_sprite[1][45][34] = 1;cactus_sprite[1][45][35] = 1;cactus_sprite[1][45][36] = 1;cactus_sprite[1][45][37] = 1;cactus_sprite[1][45][38] = 1;cactus_sprite[1][45][39] = 1;cactus_sprite[1][45][40] = 1;cactus_sprite[1][45][41] = 1;cactus_sprite[1][45][42] = 1;cactus_sprite[1][45][43] = 1;cactus_sprite[1][45][44] = 1;cactus_sprite[1][45][45] = 1;cactus_sprite[1][45][46] = 1;cactus_sprite[1][45][47] = 1;cactus_sprite[1][45][48] = 1;cactus_sprite[1][45][49] = 1;cactus_sprite[1][45][50] = 1;cactus_sprite[1][45][51] = 1;cactus_sprite[1][45][52] = 1;cactus_sprite[1][45][53] = 1;cactus_sprite[1][45][54] = 1;cactus_sprite[1][45][55] = 1;cactus_sprite[1][45][56] = 1;cactus_sprite[1][45][57] = 1;cactus_sprite[1][45][58] = 1;cactus_sprite[1][45][59] = 1;cactus_sprite[1][45][60] = 1;cactus_sprite[1][45][61] = 1;cactus_sprite[1][46][30] = 1;cactus_sprite[1][46][31] = 1;cactus_sprite[1][46][32] = 1;cactus_sprite[1][46][33] = 1;cactus_sprite[1][46][34] = 1;cactus_sprite[1][46][35] = 1;cactus_sprite[1][46][36] = 1;cactus_sprite[1][46][37] = 1;cactus_sprite[1][46][38] = 1;cactus_sprite[1][46][39] = 1;cactus_sprite[1][46][40] = 1;cactus_sprite[1][46][41] = 1;cactus_sprite[1][46][42] = 1;cactus_sprite[1][46][43] = 1;cactus_sprite[1][46][44] = 1;cactus_sprite[1][46][45] = 1;cactus_sprite[1][46][46] = 1;cactus_sprite[1][46][47] = 1;cactus_sprite[1][46][48] = 1;cactus_sprite[1][46][49] = 1;cactus_sprite[1][46][50] = 1;cactus_sprite[1][46][51] = 1;cactus_sprite[1][46][52] = 1;cactus_sprite[1][46][53] = 1;cactus_sprite[1][46][54] = 1;cactus_sprite[1][46][55] = 1;cactus_sprite[1][46][56] = 1;cactus_sprite[1][46][57] = 1;cactus_sprite[1][46][58] = 1;cactus_sprite[1][46][59] = 1;cactus_sprite[1][47][30] = 1;cactus_sprite[1][47][31] = 1;cactus_sprite[1][47][32] = 1;cactus_sprite[1][47][33] = 1;cactus_sprite[1][47][34] = 1;cactus_sprite[1][47][35] = 1;cactus_sprite[1][47][36] = 1;cactus_sprite[1][47][37] = 1;cactus_sprite[1][47][38] = 1;cactus_sprite[1][47][39] = 1;cactus_sprite[1][47][40] = 1;cactus_sprite[1][47][41] = 1;cactus_sprite[1][47][42] = 1;cactus_sprite[1][47][43] = 1;cactus_sprite[1][47][44] = 1;cactus_sprite[1][47][45] = 1;cactus_sprite[1][47][46] = 1;cactus_sprite[1][47][47] = 1;cactus_sprite[1][47][48] = 1;cactus_sprite[1][47][49] = 1;cactus_sprite[1][47][50] = 1;cactus_sprite[1][47][51] = 1;cactus_sprite[1][47][52] = 1;cactus_sprite[1][47][53] = 1;cactus_sprite[1][47][54] = 1;cactus_sprite[1][47][55] = 1;cactus_sprite[1][47][56] = 1;cactus_sprite[1][47][57] = 1;cactus_sprite[1][47][58] = 1;cactus_sprite[1][47][59] = 1;
	cactus_sprite[2][2][34] = 1;cactus_sprite[2][2][35] = 1;cactus_sprite[2][2][36] = 1;cactus_sprite[2][2][37] = 1;cactus_sprite[2][2][38] = 1;cactus_sprite[2][2][39] = 1;cactus_sprite[2][2][40] = 1;cactus_sprite[2][2][41] = 1;cactus_sprite[2][2][42] = 1;cactus_sprite[2][2][43] = 1;cactus_sprite[2][2][44] = 1;cactus_sprite[2][2][45] = 1;cactus_sprite[2][2][46] = 1;cactus_sprite[2][2][47] = 1;cactus_sprite[2][2][48] = 1;cactus_sprite[2][2][49] = 1;cactus_sprite[2][2][50] = 1;cactus_sprite[2][2][51] = 1;cactus_sprite[2][2][52] = 1;cactus_sprite[2][2][53] = 1;cactus_sprite[2][2][54] = 1;cactus_sprite[2][2][55] = 1;cactus_sprite[2][2][56] = 1;cactus_sprite[2][2][57] = 1;cactus_sprite[2][2][58] = 1;cactus_sprite[2][2][59] = 1;cactus_sprite[2][2][60] = 1;cactus_sprite[2][2][61] = 1;cactus_sprite[2][2][62] = 1;cactus_sprite[2][2][63] = 1;cactus_sprite[2][3][34] = 1;cactus_sprite[2][3][35] = 1;cactus_sprite[2][3][36] = 1;cactus_sprite[2][3][37] = 1;cactus_sprite[2][3][38] = 1;cactus_sprite[2][3][39] = 1;cactus_sprite[2][3][40] = 1;cactus_sprite[2][3][41] = 1;cactus_sprite[2][3][42] = 1;cactus_sprite[2][3][43] = 1;cactus_sprite[2][3][44] = 1;cactus_sprite[2][3][45] = 1;cactus_sprite[2][3][46] = 1;cactus_sprite[2][3][47] = 1;cactus_sprite[2][3][48] = 1;cactus_sprite[2][3][49] = 1;cactus_sprite[2][3][50] = 1;cactus_sprite[2][3][51] = 1;cactus_sprite[2][3][52] = 1;cactus_sprite[2][3][53] = 1;cactus_sprite[2][3][54] = 1;cactus_sprite[2][3][55] = 1;cactus_sprite[2][3][56] = 1;cactus_sprite[2][3][57] = 1;cactus_sprite[2][3][58] = 1;cactus_sprite[2][3][59] = 1;cactus_sprite[2][3][60] = 1;cactus_sprite[2][3][61] = 1;cactus_sprite[2][3][62] = 1;cactus_sprite[2][3][63] = 1;cactus_sprite[2][4][32] = 1;cactus_sprite[2][4][33] = 1;cactus_sprite[2][4][34] = 1;cactus_sprite[2][4][35] = 1;cactus_sprite[2][4][36] = 1;cactus_sprite[2][4][37] = 1;cactus_sprite[2][4][38] = 1;cactus_sprite[2][4][39] = 1;cactus_sprite[2][4][40] = 1;cactus_sprite[2][4][41] = 1;cactus_sprite[2][4][42] = 1;cactus_sprite[2][4][43] = 1;cactus_sprite[2][4][44] = 1;cactus_sprite[2][4][45] = 1;cactus_sprite[2][4][46] = 1;cactus_sprite[2][4][47] = 1;cactus_sprite[2][4][48] = 1;cactus_sprite[2][4][49] = 1;cactus_sprite[2][4][50] = 1;cactus_sprite[2][4][51] = 1;cactus_sprite[2][4][52] = 1;cactus_sprite[2][4][53] = 1;cactus_sprite[2][4][54] = 1;cactus_sprite[2][4][55] = 1;cactus_sprite[2][4][56] = 1;cactus_sprite[2][4][57] = 1;cactus_sprite[2][4][58] = 1;cactus_sprite[2][4][59] = 1;cactus_sprite[2][4][60] = 1;cactus_sprite[2][4][61] = 1;cactus_sprite[2][4][62] = 1;cactus_sprite[2][4][63] = 1;cactus_sprite[2][4][64] = 1;cactus_sprite[2][4][65] = 1;cactus_sprite[2][5][32] = 1;cactus_sprite[2][5][33] = 1;cactus_sprite[2][5][34] = 1;cactus_sprite[2][5][35] = 1;cactus_sprite[2][5][36] = 1;cactus_sprite[2][5][37] = 1;cactus_sprite[2][5][38] = 1;cactus_sprite[2][5][39] = 1;cactus_sprite[2][5][40] = 1;cactus_sprite[2][5][41] = 1;cactus_sprite[2][5][42] = 1;cactus_sprite[2][5][43] = 1;cactus_sprite[2][5][44] = 1;cactus_sprite[2][5][45] = 1;cactus_sprite[2][5][46] = 1;cactus_sprite[2][5][47] = 1;cactus_sprite[2][5][48] = 1;cactus_sprite[2][5][49] = 1;cactus_sprite[2][5][50] = 1;cactus_sprite[2][5][51] = 1;cactus_sprite[2][5][52] = 1;cactus_sprite[2][5][53] = 1;cactus_sprite[2][5][54] = 1;cactus_sprite[2][5][55] = 1;cactus_sprite[2][5][56] = 1;cactus_sprite[2][5][57] = 1;cactus_sprite[2][5][58] = 1;cactus_sprite[2][5][59] = 1;cactus_sprite[2][5][60] = 1;cactus_sprite[2][5][61] = 1;cactus_sprite[2][5][62] = 1;cactus_sprite[2][5][63] = 1;cactus_sprite[2][5][64] = 1;cactus_sprite[2][5][65] = 1;cactus_sprite[2][6][32] = 1;cactus_sprite[2][6][33] = 1;cactus_sprite[2][6][34] = 1;cactus_sprite[2][6][35] = 1;cactus_sprite[2][6][36] = 1;cactus_sprite[2][6][37] = 1;cactus_sprite[2][6][38] = 1;cactus_sprite[2][6][39] = 1;cactus_sprite[2][6][40] = 1;cactus_sprite[2][6][41] = 1;cactus_sprite[2][6][42] = 1;cactus_sprite[2][6][43] = 1;cactus_sprite[2][6][44] = 1;cactus_sprite[2][6][45] = 1;cactus_sprite[2][6][46] = 1;cactus_sprite[2][6][47] = 1;cactus_sprite[2][6][48] = 1;cactus_sprite[2][6][49] = 1;cactus_sprite[2][6][50] = 1;cactus_sprite[2][6][51] = 1;cactus_sprite[2][6][52] = 1;cactus_sprite[2][6][53] = 1;cactus_sprite[2][6][54] = 1;cactus_sprite[2][6][55] = 1;cactus_sprite[2][6][56] = 1;cactus_sprite[2][6][57] = 1;cactus_sprite[2][6][58] = 1;cactus_sprite[2][6][59] = 1;cactus_sprite[2][6][60] = 1;cactus_sprite[2][6][61] = 1;cactus_sprite[2][6][62] = 1;cactus_sprite[2][6][63] = 1;cactus_sprite[2][6][64] = 1;cactus_sprite[2][6][65] = 1;cactus_sprite[2][6][66] = 1;cactus_sprite[2][6][67] = 1;cactus_sprite[2][7][32] = 1;cactus_sprite[2][7][33] = 1;cactus_sprite[2][7][34] = 1;cactus_sprite[2][7][35] = 1;cactus_sprite[2][7][36] = 1;cactus_sprite[2][7][37] = 1;cactus_sprite[2][7][38] = 1;cactus_sprite[2][7][39] = 1;cactus_sprite[2][7][40] = 1;cactus_sprite[2][7][41] = 1;cactus_sprite[2][7][42] = 1;cactus_sprite[2][7][43] = 1;cactus_sprite[2][7][44] = 1;cactus_sprite[2][7][45] = 1;cactus_sprite[2][7][46] = 1;cactus_sprite[2][7][47] = 1;cactus_sprite[2][7][48] = 1;cactus_sprite[2][7][49] = 1;cactus_sprite[2][7][50] = 1;cactus_sprite[2][7][51] = 1;cactus_sprite[2][7][52] = 1;cactus_sprite[2][7][53] = 1;cactus_sprite[2][7][54] = 1;cactus_sprite[2][7][55] = 1;cactus_sprite[2][7][56] = 1;cactus_sprite[2][7][57] = 1;cactus_sprite[2][7][58] = 1;cactus_sprite[2][7][59] = 1;cactus_sprite[2][7][60] = 1;cactus_sprite[2][7][61] = 1;cactus_sprite[2][7][62] = 1;cactus_sprite[2][7][63] = 1;cactus_sprite[2][7][64] = 1;cactus_sprite[2][7][65] = 1;cactus_sprite[2][7][66] = 1;cactus_sprite[2][7][67] = 1;cactus_sprite[2][8][32] = 1;cactus_sprite[2][8][33] = 1;cactus_sprite[2][8][34] = 1;cactus_sprite[2][8][35] = 1;cactus_sprite[2][8][36] = 1;cactus_sprite[2][8][37] = 1;cactus_sprite[2][8][38] = 1;cactus_sprite[2][8][39] = 1;cactus_sprite[2][8][40] = 1;cactus_sprite[2][8][41] = 1;cactus_sprite[2][8][42] = 1;cactus_sprite[2][8][43] = 1;cactus_sprite[2][8][44] = 1;cactus_sprite[2][8][45] = 1;cactus_sprite[2][8][46] = 1;cactus_sprite[2][8][47] = 1;cactus_sprite[2][8][48] = 1;cactus_sprite[2][8][49] = 1;cactus_sprite[2][8][50] = 1;cactus_sprite[2][8][51] = 1;cactus_sprite[2][8][52] = 1;cactus_sprite[2][8][53] = 1;cactus_sprite[2][8][54] = 1;cactus_sprite[2][8][55] = 1;cactus_sprite[2][8][56] = 1;cactus_sprite[2][8][57] = 1;cactus_sprite[2][8][58] = 1;cactus_sprite[2][8][59] = 1;cactus_sprite[2][8][60] = 1;cactus_sprite[2][8][61] = 1;cactus_sprite[2][8][62] = 1;cactus_sprite[2][8][63] = 1;cactus_sprite[2][8][64] = 1;cactus_sprite[2][8][65] = 1;cactus_sprite[2][8][66] = 1;cactus_sprite[2][8][67] = 1;cactus_sprite[2][8][68] = 1;cactus_sprite[2][8][69] = 1;cactus_sprite[2][9][32] = 1;cactus_sprite[2][9][33] = 1;cactus_sprite[2][9][34] = 1;cactus_sprite[2][9][35] = 1;cactus_sprite[2][9][36] = 1;cactus_sprite[2][9][37] = 1;cactus_sprite[2][9][38] = 1;cactus_sprite[2][9][39] = 1;cactus_sprite[2][9][40] = 1;cactus_sprite[2][9][41] = 1;cactus_sprite[2][9][42] = 1;cactus_sprite[2][9][43] = 1;cactus_sprite[2][9][44] = 1;cactus_sprite[2][9][45] = 1;cactus_sprite[2][9][46] = 1;cactus_sprite[2][9][47] = 1;cactus_sprite[2][9][48] = 1;cactus_sprite[2][9][49] = 1;cactus_sprite[2][9][50] = 1;cactus_sprite[2][9][51] = 1;cactus_sprite[2][9][52] = 1;cactus_sprite[2][9][53] = 1;cactus_sprite[2][9][54] = 1;cactus_sprite[2][9][55] = 1;cactus_sprite[2][9][56] = 1;cactus_sprite[2][9][57] = 1;cactus_sprite[2][9][58] = 1;cactus_sprite[2][9][59] = 1;cactus_sprite[2][9][60] = 1;cactus_sprite[2][9][61] = 1;cactus_sprite[2][9][62] = 1;cactus_sprite[2][9][63] = 1;cactus_sprite[2][9][64] = 1;cactus_sprite[2][9][65] = 1;cactus_sprite[2][9][66] = 1;cactus_sprite[2][9][67] = 1;cactus_sprite[2][9][68] = 1;cactus_sprite[2][9][69] = 1;cactus_sprite[2][10][34] = 1;cactus_sprite[2][10][35] = 1;cactus_sprite[2][10][36] = 1;cactus_sprite[2][10][37] = 1;cactus_sprite[2][10][38] = 1;cactus_sprite[2][10][39] = 1;cactus_sprite[2][10][40] = 1;cactus_sprite[2][10][41] = 1;cactus_sprite[2][10][42] = 1;cactus_sprite[2][10][43] = 1;cactus_sprite[2][10][44] = 1;cactus_sprite[2][10][45] = 1;cactus_sprite[2][10][46] = 1;cactus_sprite[2][10][47] = 1;cactus_sprite[2][10][48] = 1;cactus_sprite[2][10][49] = 1;cactus_sprite[2][10][50] = 1;cactus_sprite[2][10][51] = 1;cactus_sprite[2][10][52] = 1;cactus_sprite[2][10][53] = 1;cactus_sprite[2][10][54] = 1;cactus_sprite[2][10][55] = 1;cactus_sprite[2][10][56] = 1;cactus_sprite[2][10][57] = 1;cactus_sprite[2][10][58] = 1;cactus_sprite[2][10][59] = 1;cactus_sprite[2][10][60] = 1;cactus_sprite[2][10][61] = 1;cactus_sprite[2][10][62] = 1;cactus_sprite[2][10][63] = 1;cactus_sprite[2][10][64] = 1;cactus_sprite[2][10][65] = 1;cactus_sprite[2][10][66] = 1;cactus_sprite[2][10][67] = 1;cactus_sprite[2][10][68] = 1;cactus_sprite[2][10][69] = 1;cactus_sprite[2][11][34] = 1;cactus_sprite[2][11][35] = 1;cactus_sprite[2][11][36] = 1;cactus_sprite[2][11][37] = 1;cactus_sprite[2][11][38] = 1;cactus_sprite[2][11][39] = 1;cactus_sprite[2][11][40] = 1;cactus_sprite[2][11][41] = 1;cactus_sprite[2][11][42] = 1;cactus_sprite[2][11][43] = 1;cactus_sprite[2][11][44] = 1;cactus_sprite[2][11][45] = 1;cactus_sprite[2][11][46] = 1;cactus_sprite[2][11][47] = 1;cactus_sprite[2][11][48] = 1;cactus_sprite[2][11][49] = 1;cactus_sprite[2][11][50] = 1;cactus_sprite[2][11][51] = 1;cactus_sprite[2][11][52] = 1;cactus_sprite[2][11][53] = 1;cactus_sprite[2][11][54] = 1;cactus_sprite[2][11][55] = 1;cactus_sprite[2][11][56] = 1;cactus_sprite[2][11][57] = 1;cactus_sprite[2][11][58] = 1;cactus_sprite[2][11][59] = 1;cactus_sprite[2][11][60] = 1;cactus_sprite[2][11][61] = 1;cactus_sprite[2][11][62] = 1;cactus_sprite[2][11][63] = 1;cactus_sprite[2][11][64] = 1;cactus_sprite[2][11][65] = 1;cactus_sprite[2][11][66] = 1;cactus_sprite[2][11][67] = 1;cactus_sprite[2][11][68] = 1;cactus_sprite[2][11][69] = 1;cactus_sprite[2][12][60] = 1;cactus_sprite[2][12][61] = 1;cactus_sprite[2][12][62] = 1;cactus_sprite[2][12][63] = 1;cactus_sprite[2][12][64] = 1;cactus_sprite[2][12][65] = 1;cactus_sprite[2][12][66] = 1;cactus_sprite[2][12][67] = 1;cactus_sprite[2][12][68] = 1;cactus_sprite[2][12][69] = 1;cactus_sprite[2][13][60] = 1;cactus_sprite[2][13][61] = 1;cactus_sprite[2][13][62] = 1;cactus_sprite[2][13][63] = 1;cactus_sprite[2][13][64] = 1;cactus_sprite[2][13][65] = 1;cactus_sprite[2][13][66] = 1;cactus_sprite[2][13][67] = 1;cactus_sprite[2][13][68] = 1;cactus_sprite[2][13][69] = 1;cactus_sprite[2][14][60] = 1;cactus_sprite[2][14][61] = 1;cactus_sprite[2][14][62] = 1;cactus_sprite[2][14][63] = 1;cactus_sprite[2][14][64] = 1;cactus_sprite[2][14][65] = 1;cactus_sprite[2][14][66] = 1;cactus_sprite[2][14][67] = 1;cactus_sprite[2][14][68] = 1;cactus_sprite[2][14][69] = 1;cactus_sprite[2][15][60] = 1;cactus_sprite[2][15][61] = 1;cactus_sprite[2][15][62] = 1;cactus_sprite[2][15][63] = 1;cactus_sprite[2][15][64] = 1;cactus_sprite[2][15][65] = 1;cactus_sprite[2][15][66] = 1;cactus_sprite[2][15][67] = 1;cactus_sprite[2][15][68] = 1;cactus_sprite[2][15][69] = 1;cactus_sprite[2][16][60] = 1;cactus_sprite[2][16][61] = 1;cactus_sprite[2][16][62] = 1;cactus_sprite[2][16][63] = 1;cactus_sprite[2][16][64] = 1;cactus_sprite[2][16][65] = 1;cactus_sprite[2][16][66] = 1;cactus_sprite[2][16][67] = 1;cactus_sprite[2][16][68] = 1;cactus_sprite[2][16][69] = 1;cactus_sprite[2][17][60] = 1;cactus_sprite[2][17][61] = 1;cactus_sprite[2][17][62] = 1;cactus_sprite[2][17][63] = 1;cactus_sprite[2][17][64] = 1;cactus_sprite[2][17][65] = 1;cactus_sprite[2][17][66] = 1;cactus_sprite[2][17][67] = 1;cactus_sprite[2][17][68] = 1;cactus_sprite[2][17][69] = 1;cactus_sprite[2][18][10] = 1;cactus_sprite[2][18][11] = 1;cactus_sprite[2][18][12] = 1;cactus_sprite[2][18][13] = 1;cactus_sprite[2][18][14] = 1;cactus_sprite[2][18][15] = 1;cactus_sprite[2][18][16] = 1;cactus_sprite[2][18][17] = 1;cactus_sprite[2][18][18] = 1;cactus_sprite[2][18][19] = 1;cactus_sprite[2][18][20] = 1;cactus_sprite[2][18][21] = 1;cactus_sprite[2][18][22] = 1;cactus_sprite[2][18][23] = 1;cactus_sprite[2][18][24] = 1;cactus_sprite[2][18][25] = 1;cactus_sprite[2][18][26] = 1;cactus_sprite[2][18][27] = 1;cactus_sprite[2][18][28] = 1;cactus_sprite[2][18][29] = 1;cactus_sprite[2][18][30] = 1;cactus_sprite[2][18][31] = 1;cactus_sprite[2][18][32] = 1;cactus_sprite[2][18][33] = 1;cactus_sprite[2][18][34] = 1;cactus_sprite[2][18][35] = 1;cactus_sprite[2][18][36] = 1;cactus_sprite[2][18][37] = 1;cactus_sprite[2][18][38] = 1;cactus_sprite[2][18][39] = 1;cactus_sprite[2][18][40] = 1;cactus_sprite[2][18][41] = 1;cactus_sprite[2][18][42] = 1;cactus_sprite[2][18][43] = 1;cactus_sprite[2][18][44] = 1;cactus_sprite[2][18][45] = 1;cactus_sprite[2][18][46] = 1;cactus_sprite[2][18][47] = 1;cactus_sprite[2][18][48] = 1;cactus_sprite[2][18][49] = 1;cactus_sprite[2][18][50] = 1;cactus_sprite[2][18][51] = 1;cactus_sprite[2][18][52] = 1;cactus_sprite[2][18][53] = 1;cactus_sprite[2][18][54] = 1;cactus_sprite[2][18][55] = 1;cactus_sprite[2][18][56] = 1;cactus_sprite[2][18][57] = 1;cactus_sprite[2][18][58] = 1;cactus_sprite[2][18][59] = 1;cactus_sprite[2][18][60] = 1;cactus_sprite[2][18][61] = 1;cactus_sprite[2][18][62] = 1;cactus_sprite[2][18][63] = 1;cactus_sprite[2][18][64] = 1;cactus_sprite[2][18][65] = 1;cactus_sprite[2][18][66] = 1;cactus_sprite[2][18][67] = 1;cactus_sprite[2][18][68] = 1;cactus_sprite[2][18][69] = 1;cactus_sprite[2][18][70] = 1;cactus_sprite[2][18][71] = 1;cactus_sprite[2][18][72] = 1;cactus_sprite[2][18][73] = 1;cactus_sprite[2][18][74] = 1;cactus_sprite[2][18][75] = 1;cactus_sprite[2][18][76] = 1;cactus_sprite[2][18][77] = 1;cactus_sprite[2][18][78] = 1;cactus_sprite[2][18][79] = 1;cactus_sprite[2][18][80] = 1;cactus_sprite[2][18][81] = 1;cactus_sprite[2][18][82] = 1;cactus_sprite[2][18][83] = 1;cactus_sprite[2][18][84] = 1;cactus_sprite[2][18][85] = 1;cactus_sprite[2][18][86] = 1;cactus_sprite[2][18][87] = 1;cactus_sprite[2][18][88] = 1;cactus_sprite[2][18][89] = 1;cactus_sprite[2][18][90] = 1;cactus_sprite[2][18][91] = 1;cactus_sprite[2][18][92] = 1;cactus_sprite[2][18][93] = 1;cactus_sprite[2][18][94] = 1;cactus_sprite[2][18][95] = 1;cactus_sprite[2][18][96] = 1;cactus_sprite[2][18][97] = 1;cactus_sprite[2][18][98] = 1;cactus_sprite[2][18][99] = 1;cactus_sprite[2][19][10] = 1;cactus_sprite[2][19][11] = 1;cactus_sprite[2][19][12] = 1;cactus_sprite[2][19][13] = 1;cactus_sprite[2][19][14] = 1;cactus_sprite[2][19][15] = 1;cactus_sprite[2][19][16] = 1;cactus_sprite[2][19][17] = 1;cactus_sprite[2][19][18] = 1;cactus_sprite[2][19][19] = 1;cactus_sprite[2][19][20] = 1;cactus_sprite[2][19][21] = 1;cactus_sprite[2][19][22] = 1;cactus_sprite[2][19][23] = 1;cactus_sprite[2][19][24] = 1;cactus_sprite[2][19][25] = 1;cactus_sprite[2][19][26] = 1;cactus_sprite[2][19][27] = 1;cactus_sprite[2][19][28] = 1;cactus_sprite[2][19][29] = 1;cactus_sprite[2][19][30] = 1;cactus_sprite[2][19][31] = 1;cactus_sprite[2][19][32] = 1;cactus_sprite[2][19][33] = 1;cactus_sprite[2][19][34] = 1;cactus_sprite[2][19][35] = 1;cactus_sprite[2][19][36] = 1;cactus_sprite[2][19][37] = 1;cactus_sprite[2][19][38] = 1;cactus_sprite[2][19][39] = 1;cactus_sprite[2][19][40] = 1;cactus_sprite[2][19][41] = 1;cactus_sprite[2][19][42] = 1;cactus_sprite[2][19][43] = 1;cactus_sprite[2][19][44] = 1;cactus_sprite[2][19][45] = 1;cactus_sprite[2][19][46] = 1;cactus_sprite[2][19][47] = 1;cactus_sprite[2][19][48] = 1;cactus_sprite[2][19][49] = 1;cactus_sprite[2][19][50] = 1;cactus_sprite[2][19][51] = 1;cactus_sprite[2][19][52] = 1;cactus_sprite[2][19][53] = 1;cactus_sprite[2][19][54] = 1;cactus_sprite[2][19][55] = 1;cactus_sprite[2][19][56] = 1;cactus_sprite[2][19][57] = 1;cactus_sprite[2][19][58] = 1;cactus_sprite[2][19][59] = 1;cactus_sprite[2][19][60] = 1;cactus_sprite[2][19][61] = 1;cactus_sprite[2][19][62] = 1;cactus_sprite[2][19][63] = 1;cactus_sprite[2][19][64] = 1;cactus_sprite[2][19][65] = 1;cactus_sprite[2][19][66] = 1;cactus_sprite[2][19][67] = 1;cactus_sprite[2][19][68] = 1;cactus_sprite[2][19][69] = 1;cactus_sprite[2][19][70] = 1;cactus_sprite[2][19][71] = 1;cactus_sprite[2][19][72] = 1;cactus_sprite[2][19][73] = 1;cactus_sprite[2][19][74] = 1;cactus_sprite[2][19][75] = 1;cactus_sprite[2][19][76] = 1;cactus_sprite[2][19][77] = 1;cactus_sprite[2][19][78] = 1;cactus_sprite[2][19][79] = 1;cactus_sprite[2][19][80] = 1;cactus_sprite[2][19][81] = 1;cactus_sprite[2][19][82] = 1;cactus_sprite[2][19][83] = 1;cactus_sprite[2][19][84] = 1;cactus_sprite[2][19][85] = 1;cactus_sprite[2][19][86] = 1;cactus_sprite[2][19][87] = 1;cactus_sprite[2][19][88] = 1;cactus_sprite[2][19][89] = 1;cactus_sprite[2][19][90] = 1;cactus_sprite[2][19][91] = 1;cactus_sprite[2][19][92] = 1;cactus_sprite[2][19][93] = 1;cactus_sprite[2][19][94] = 1;cactus_sprite[2][19][95] = 1;cactus_sprite[2][19][96] = 1;cactus_sprite[2][19][97] = 1;cactus_sprite[2][19][98] = 1;cactus_sprite[2][19][99] = 1;cactus_sprite[2][20][8] = 1;cactus_sprite[2][20][9] = 1;cactus_sprite[2][20][10] = 1;cactus_sprite[2][20][11] = 1;cactus_sprite[2][20][12] = 1;cactus_sprite[2][20][13] = 1;cactus_sprite[2][20][14] = 1;cactus_sprite[2][20][15] = 1;cactus_sprite[2][20][16] = 1;cactus_sprite[2][20][17] = 1;cactus_sprite[2][20][18] = 1;cactus_sprite[2][20][19] = 1;cactus_sprite[2][20][20] = 1;cactus_sprite[2][20][21] = 1;cactus_sprite[2][20][22] = 1;cactus_sprite[2][20][23] = 1;cactus_sprite[2][20][24] = 1;cactus_sprite[2][20][25] = 1;cactus_sprite[2][20][26] = 1;cactus_sprite[2][20][27] = 1;cactus_sprite[2][20][28] = 1;cactus_sprite[2][20][29] = 1;cactus_sprite[2][20][30] = 1;cactus_sprite[2][20][31] = 1;cactus_sprite[2][20][32] = 1;cactus_sprite[2][20][33] = 1;cactus_sprite[2][20][34] = 1;cactus_sprite[2][20][35] = 1;cactus_sprite[2][20][36] = 1;cactus_sprite[2][20][37] = 1;cactus_sprite[2][20][38] = 1;cactus_sprite[2][20][39] = 1;cactus_sprite[2][20][40] = 1;cactus_sprite[2][20][41] = 1;cactus_sprite[2][20][42] = 1;cactus_sprite[2][20][43] = 1;cactus_sprite[2][20][44] = 1;cactus_sprite[2][20][45] = 1;cactus_sprite[2][20][46] = 1;cactus_sprite[2][20][47] = 1;cactus_sprite[2][20][48] = 1;cactus_sprite[2][20][49] = 1;cactus_sprite[2][20][50] = 1;cactus_sprite[2][20][51] = 1;cactus_sprite[2][20][52] = 1;cactus_sprite[2][20][53] = 1;cactus_sprite[2][20][54] = 1;cactus_sprite[2][20][55] = 1;cactus_sprite[2][20][56] = 1;cactus_sprite[2][20][57] = 1;cactus_sprite[2][20][58] = 1;cactus_sprite[2][20][59] = 1;cactus_sprite[2][20][60] = 1;cactus_sprite[2][20][61] = 1;cactus_sprite[2][20][62] = 1;cactus_sprite[2][20][63] = 1;cactus_sprite[2][20][64] = 1;cactus_sprite[2][20][65] = 1;cactus_sprite[2][20][66] = 1;cactus_sprite[2][20][67] = 1;cactus_sprite[2][20][68] = 1;cactus_sprite[2][20][69] = 1;cactus_sprite[2][20][70] = 1;cactus_sprite[2][20][71] = 1;cactus_sprite[2][20][72] = 1;cactus_sprite[2][20][73] = 1;cactus_sprite[2][20][74] = 1;cactus_sprite[2][20][75] = 1;cactus_sprite[2][20][76] = 1;cactus_sprite[2][20][77] = 1;cactus_sprite[2][20][78] = 1;cactus_sprite[2][20][79] = 1;cactus_sprite[2][20][80] = 1;cactus_sprite[2][20][81] = 1;cactus_sprite[2][20][82] = 1;cactus_sprite[2][20][83] = 1;cactus_sprite[2][20][84] = 1;cactus_sprite[2][20][85] = 1;cactus_sprite[2][20][86] = 1;cactus_sprite[2][20][87] = 1;cactus_sprite[2][20][88] = 1;cactus_sprite[2][20][89] = 1;cactus_sprite[2][20][90] = 1;cactus_sprite[2][20][91] = 1;cactus_sprite[2][20][92] = 1;cactus_sprite[2][20][93] = 1;cactus_sprite[2][20][94] = 1;cactus_sprite[2][20][95] = 1;cactus_sprite[2][20][96] = 1;cactus_sprite[2][20][97] = 1;cactus_sprite[2][20][98] = 1;cactus_sprite[2][20][99] = 1;cactus_sprite[2][21][8] = 1;cactus_sprite[2][21][9] = 1;cactus_sprite[2][21][10] = 1;cactus_sprite[2][21][11] = 1;cactus_sprite[2][21][12] = 1;cactus_sprite[2][21][13] = 1;cactus_sprite[2][21][14] = 1;cactus_sprite[2][21][15] = 1;cactus_sprite[2][21][16] = 1;cactus_sprite[2][21][17] = 1;cactus_sprite[2][21][18] = 1;cactus_sprite[2][21][19] = 1;cactus_sprite[2][21][20] = 1;cactus_sprite[2][21][21] = 1;cactus_sprite[2][21][22] = 1;cactus_sprite[2][21][23] = 1;cactus_sprite[2][21][24] = 1;cactus_sprite[2][21][25] = 1;cactus_sprite[2][21][26] = 1;cactus_sprite[2][21][27] = 1;cactus_sprite[2][21][28] = 1;cactus_sprite[2][21][29] = 1;cactus_sprite[2][21][30] = 1;cactus_sprite[2][21][31] = 1;cactus_sprite[2][21][32] = 1;cactus_sprite[2][21][33] = 1;cactus_sprite[2][21][34] = 1;cactus_sprite[2][21][35] = 1;cactus_sprite[2][21][36] = 1;cactus_sprite[2][21][37] = 1;cactus_sprite[2][21][38] = 1;cactus_sprite[2][21][39] = 1;cactus_sprite[2][21][40] = 1;cactus_sprite[2][21][41] = 1;cactus_sprite[2][21][42] = 1;cactus_sprite[2][21][43] = 1;cactus_sprite[2][21][44] = 1;cactus_sprite[2][21][45] = 1;cactus_sprite[2][21][46] = 1;cactus_sprite[2][21][47] = 1;cactus_sprite[2][21][48] = 1;cactus_sprite[2][21][49] = 1;cactus_sprite[2][21][50] = 1;cactus_sprite[2][21][51] = 1;cactus_sprite[2][21][52] = 1;cactus_sprite[2][21][53] = 1;cactus_sprite[2][21][54] = 1;cactus_sprite[2][21][55] = 1;cactus_sprite[2][21][56] = 1;cactus_sprite[2][21][57] = 1;cactus_sprite[2][21][58] = 1;cactus_sprite[2][21][59] = 1;cactus_sprite[2][21][60] = 1;cactus_sprite[2][21][61] = 1;cactus_sprite[2][21][62] = 1;cactus_sprite[2][21][63] = 1;cactus_sprite[2][21][64] = 1;cactus_sprite[2][21][65] = 1;cactus_sprite[2][21][66] = 1;cactus_sprite[2][21][67] = 1;cactus_sprite[2][21][68] = 1;cactus_sprite[2][21][69] = 1;cactus_sprite[2][21][70] = 1;cactus_sprite[2][21][71] = 1;cactus_sprite[2][21][72] = 1;cactus_sprite[2][21][73] = 1;cactus_sprite[2][21][74] = 1;cactus_sprite[2][21][75] = 1;cactus_sprite[2][21][76] = 1;cactus_sprite[2][21][77] = 1;cactus_sprite[2][21][78] = 1;cactus_sprite[2][21][79] = 1;cactus_sprite[2][21][80] = 1;cactus_sprite[2][21][81] = 1;cactus_sprite[2][21][82] = 1;cactus_sprite[2][21][83] = 1;cactus_sprite[2][21][84] = 1;cactus_sprite[2][21][85] = 1;cactus_sprite[2][21][86] = 1;cactus_sprite[2][21][87] = 1;cactus_sprite[2][21][88] = 1;cactus_sprite[2][21][89] = 1;cactus_sprite[2][21][90] = 1;cactus_sprite[2][21][91] = 1;cactus_sprite[2][21][92] = 1;cactus_sprite[2][21][93] = 1;cactus_sprite[2][21][94] = 1;cactus_sprite[2][21][95] = 1;cactus_sprite[2][21][96] = 1;cactus_sprite[2][21][97] = 1;cactus_sprite[2][21][98] = 1;cactus_sprite[2][21][99] = 1;cactus_sprite[2][22][8] = 1;cactus_sprite[2][22][9] = 1;cactus_sprite[2][22][10] = 1;cactus_sprite[2][22][11] = 1;cactus_sprite[2][22][12] = 1;cactus_sprite[2][22][13] = 1;cactus_sprite[2][22][14] = 1;cactus_sprite[2][22][15] = 1;cactus_sprite[2][22][16] = 1;cactus_sprite[2][22][17] = 1;cactus_sprite[2][22][18] = 1;cactus_sprite[2][22][19] = 1;cactus_sprite[2][22][20] = 1;cactus_sprite[2][22][21] = 1;cactus_sprite[2][22][22] = 1;cactus_sprite[2][22][23] = 1;cactus_sprite[2][22][24] = 1;cactus_sprite[2][22][25] = 1;cactus_sprite[2][22][26] = 1;cactus_sprite[2][22][27] = 1;cactus_sprite[2][22][28] = 1;cactus_sprite[2][22][29] = 1;cactus_sprite[2][22][30] = 1;cactus_sprite[2][22][31] = 1;cactus_sprite[2][22][32] = 1;cactus_sprite[2][22][33] = 1;cactus_sprite[2][22][34] = 1;cactus_sprite[2][22][35] = 1;cactus_sprite[2][22][36] = 1;cactus_sprite[2][22][37] = 1;cactus_sprite[2][22][38] = 1;cactus_sprite[2][22][39] = 1;cactus_sprite[2][22][40] = 1;cactus_sprite[2][22][41] = 1;cactus_sprite[2][22][42] = 1;cactus_sprite[2][22][43] = 1;cactus_sprite[2][22][44] = 1;cactus_sprite[2][22][45] = 1;cactus_sprite[2][22][46] = 1;cactus_sprite[2][22][47] = 1;cactus_sprite[2][22][48] = 1;cactus_sprite[2][22][49] = 1;cactus_sprite[2][22][50] = 1;cactus_sprite[2][22][51] = 1;cactus_sprite[2][22][52] = 1;cactus_sprite[2][22][53] = 1;cactus_sprite[2][22][54] = 1;cactus_sprite[2][22][55] = 1;cactus_sprite[2][22][56] = 1;cactus_sprite[2][22][57] = 1;cactus_sprite[2][22][58] = 1;cactus_sprite[2][22][59] = 1;cactus_sprite[2][22][60] = 1;cactus_sprite[2][22][61] = 1;cactus_sprite[2][22][62] = 1;cactus_sprite[2][22][63] = 1;cactus_sprite[2][22][64] = 1;cactus_sprite[2][22][65] = 1;cactus_sprite[2][22][66] = 1;cactus_sprite[2][22][67] = 1;cactus_sprite[2][22][68] = 1;cactus_sprite[2][22][69] = 1;cactus_sprite[2][22][70] = 1;cactus_sprite[2][22][71] = 1;cactus_sprite[2][22][72] = 1;cactus_sprite[2][22][73] = 1;cactus_sprite[2][22][74] = 1;cactus_sprite[2][22][75] = 1;cactus_sprite[2][22][76] = 1;cactus_sprite[2][22][77] = 1;cactus_sprite[2][22][78] = 1;cactus_sprite[2][22][79] = 1;cactus_sprite[2][22][80] = 1;cactus_sprite[2][22][81] = 1;cactus_sprite[2][22][82] = 1;cactus_sprite[2][22][83] = 1;cactus_sprite[2][22][84] = 1;cactus_sprite[2][22][85] = 1;cactus_sprite[2][22][86] = 1;cactus_sprite[2][22][87] = 1;cactus_sprite[2][22][88] = 1;cactus_sprite[2][22][89] = 1;cactus_sprite[2][22][90] = 1;cactus_sprite[2][22][91] = 1;cactus_sprite[2][22][92] = 1;cactus_sprite[2][22][93] = 1;cactus_sprite[2][22][94] = 1;cactus_sprite[2][22][95] = 1;cactus_sprite[2][22][96] = 1;cactus_sprite[2][22][97] = 1;cactus_sprite[2][22][98] = 1;cactus_sprite[2][22][99] = 1;cactus_sprite[2][23][8] = 1;cactus_sprite[2][23][9] = 1;cactus_sprite[2][23][10] = 1;cactus_sprite[2][23][11] = 1;cactus_sprite[2][23][12] = 1;cactus_sprite[2][23][13] = 1;cactus_sprite[2][23][14] = 1;cactus_sprite[2][23][15] = 1;cactus_sprite[2][23][16] = 1;cactus_sprite[2][23][17] = 1;cactus_sprite[2][23][18] = 1;cactus_sprite[2][23][19] = 1;cactus_sprite[2][23][20] = 1;cactus_sprite[2][23][21] = 1;cactus_sprite[2][23][22] = 1;cactus_sprite[2][23][23] = 1;cactus_sprite[2][23][24] = 1;cactus_sprite[2][23][25] = 1;cactus_sprite[2][23][26] = 1;cactus_sprite[2][23][27] = 1;cactus_sprite[2][23][28] = 1;cactus_sprite[2][23][29] = 1;cactus_sprite[2][23][30] = 1;cactus_sprite[2][23][31] = 1;cactus_sprite[2][23][32] = 1;cactus_sprite[2][23][33] = 1;cactus_sprite[2][23][34] = 1;cactus_sprite[2][23][35] = 1;cactus_sprite[2][23][36] = 1;cactus_sprite[2][23][37] = 1;cactus_sprite[2][23][38] = 1;cactus_sprite[2][23][39] = 1;cactus_sprite[2][23][40] = 1;cactus_sprite[2][23][41] = 1;cactus_sprite[2][23][42] = 1;cactus_sprite[2][23][43] = 1;cactus_sprite[2][23][44] = 1;cactus_sprite[2][23][45] = 1;cactus_sprite[2][23][46] = 1;cactus_sprite[2][23][47] = 1;cactus_sprite[2][23][48] = 1;cactus_sprite[2][23][49] = 1;cactus_sprite[2][23][50] = 1;cactus_sprite[2][23][51] = 1;cactus_sprite[2][23][52] = 1;cactus_sprite[2][23][53] = 1;cactus_sprite[2][23][54] = 1;cactus_sprite[2][23][55] = 1;cactus_sprite[2][23][56] = 1;cactus_sprite[2][23][57] = 1;cactus_sprite[2][23][58] = 1;cactus_sprite[2][23][59] = 1;cactus_sprite[2][23][60] = 1;cactus_sprite[2][23][61] = 1;cactus_sprite[2][23][62] = 1;cactus_sprite[2][23][63] = 1;cactus_sprite[2][23][64] = 1;cactus_sprite[2][23][65] = 1;cactus_sprite[2][23][66] = 1;cactus_sprite[2][23][67] = 1;cactus_sprite[2][23][68] = 1;cactus_sprite[2][23][69] = 1;cactus_sprite[2][23][70] = 1;cactus_sprite[2][23][71] = 1;cactus_sprite[2][23][72] = 1;cactus_sprite[2][23][73] = 1;cactus_sprite[2][23][74] = 1;cactus_sprite[2][23][75] = 1;cactus_sprite[2][23][76] = 1;cactus_sprite[2][23][77] = 1;cactus_sprite[2][23][78] = 1;cactus_sprite[2][23][79] = 1;cactus_sprite[2][23][80] = 1;cactus_sprite[2][23][81] = 1;cactus_sprite[2][23][82] = 1;cactus_sprite[2][23][83] = 1;cactus_sprite[2][23][84] = 1;cactus_sprite[2][23][85] = 1;cactus_sprite[2][23][86] = 1;cactus_sprite[2][23][87] = 1;cactus_sprite[2][23][88] = 1;cactus_sprite[2][23][89] = 1;cactus_sprite[2][23][90] = 1;cactus_sprite[2][23][91] = 1;cactus_sprite[2][23][92] = 1;cactus_sprite[2][23][93] = 1;cactus_sprite[2][23][94] = 1;cactus_sprite[2][23][95] = 1;cactus_sprite[2][23][96] = 1;cactus_sprite[2][23][97] = 1;cactus_sprite[2][23][98] = 1;cactus_sprite[2][23][99] = 1;cactus_sprite[2][24][8] = 1;cactus_sprite[2][24][9] = 1;cactus_sprite[2][24][10] = 1;cactus_sprite[2][24][11] = 1;cactus_sprite[2][24][12] = 1;cactus_sprite[2][24][13] = 1;cactus_sprite[2][24][14] = 1;cactus_sprite[2][24][15] = 1;cactus_sprite[2][24][16] = 1;cactus_sprite[2][24][17] = 1;cactus_sprite[2][24][18] = 1;cactus_sprite[2][24][19] = 1;cactus_sprite[2][24][20] = 1;cactus_sprite[2][24][21] = 1;cactus_sprite[2][24][22] = 1;cactus_sprite[2][24][23] = 1;cactus_sprite[2][24][24] = 1;cactus_sprite[2][24][25] = 1;cactus_sprite[2][24][26] = 1;cactus_sprite[2][24][27] = 1;cactus_sprite[2][24][28] = 1;cactus_sprite[2][24][29] = 1;cactus_sprite[2][24][30] = 1;cactus_sprite[2][24][31] = 1;cactus_sprite[2][24][32] = 1;cactus_sprite[2][24][33] = 1;cactus_sprite[2][24][34] = 1;cactus_sprite[2][24][35] = 1;cactus_sprite[2][24][36] = 1;cactus_sprite[2][24][37] = 1;cactus_sprite[2][24][38] = 1;cactus_sprite[2][24][39] = 1;cactus_sprite[2][24][40] = 1;cactus_sprite[2][24][41] = 1;cactus_sprite[2][24][42] = 1;cactus_sprite[2][24][43] = 1;cactus_sprite[2][24][44] = 1;cactus_sprite[2][24][45] = 1;cactus_sprite[2][24][46] = 1;cactus_sprite[2][24][47] = 1;cactus_sprite[2][24][48] = 1;cactus_sprite[2][24][49] = 1;cactus_sprite[2][24][50] = 1;cactus_sprite[2][24][51] = 1;cactus_sprite[2][24][52] = 1;cactus_sprite[2][24][53] = 1;cactus_sprite[2][24][54] = 1;cactus_sprite[2][24][55] = 1;cactus_sprite[2][24][56] = 1;cactus_sprite[2][24][57] = 1;cactus_sprite[2][24][58] = 1;cactus_sprite[2][24][59] = 1;cactus_sprite[2][24][60] = 1;cactus_sprite[2][24][61] = 1;cactus_sprite[2][24][62] = 1;cactus_sprite[2][24][63] = 1;cactus_sprite[2][24][64] = 1;cactus_sprite[2][24][65] = 1;cactus_sprite[2][24][66] = 1;cactus_sprite[2][24][67] = 1;cactus_sprite[2][24][68] = 1;cactus_sprite[2][24][69] = 1;cactus_sprite[2][24][70] = 1;cactus_sprite[2][24][71] = 1;cactus_sprite[2][24][72] = 1;cactus_sprite[2][24][73] = 1;cactus_sprite[2][24][74] = 1;cactus_sprite[2][24][75] = 1;cactus_sprite[2][24][76] = 1;cactus_sprite[2][24][77] = 1;cactus_sprite[2][24][78] = 1;cactus_sprite[2][24][79] = 1;cactus_sprite[2][24][80] = 1;cactus_sprite[2][24][81] = 1;cactus_sprite[2][24][82] = 1;cactus_sprite[2][24][83] = 1;cactus_sprite[2][24][84] = 1;cactus_sprite[2][24][85] = 1;cactus_sprite[2][24][86] = 1;cactus_sprite[2][24][87] = 1;cactus_sprite[2][24][88] = 1;cactus_sprite[2][24][89] = 1;cactus_sprite[2][24][90] = 1;cactus_sprite[2][24][91] = 1;cactus_sprite[2][24][92] = 1;cactus_sprite[2][24][93] = 1;cactus_sprite[2][24][94] = 1;cactus_sprite[2][24][95] = 1;cactus_sprite[2][24][96] = 1;cactus_sprite[2][24][97] = 1;cactus_sprite[2][24][98] = 1;cactus_sprite[2][24][99] = 1;cactus_sprite[2][25][8] = 1;cactus_sprite[2][25][9] = 1;cactus_sprite[2][25][10] = 1;cactus_sprite[2][25][11] = 1;cactus_sprite[2][25][12] = 1;cactus_sprite[2][25][13] = 1;cactus_sprite[2][25][14] = 1;cactus_sprite[2][25][15] = 1;cactus_sprite[2][25][16] = 1;cactus_sprite[2][25][17] = 1;cactus_sprite[2][25][18] = 1;cactus_sprite[2][25][19] = 1;cactus_sprite[2][25][20] = 1;cactus_sprite[2][25][21] = 1;cactus_sprite[2][25][22] = 1;cactus_sprite[2][25][23] = 1;cactus_sprite[2][25][24] = 1;cactus_sprite[2][25][25] = 1;cactus_sprite[2][25][26] = 1;cactus_sprite[2][25][27] = 1;cactus_sprite[2][25][28] = 1;cactus_sprite[2][25][29] = 1;cactus_sprite[2][25][30] = 1;cactus_sprite[2][25][31] = 1;cactus_sprite[2][25][32] = 1;cactus_sprite[2][25][33] = 1;cactus_sprite[2][25][34] = 1;cactus_sprite[2][25][35] = 1;cactus_sprite[2][25][36] = 1;cactus_sprite[2][25][37] = 1;cactus_sprite[2][25][38] = 1;cactus_sprite[2][25][39] = 1;cactus_sprite[2][25][40] = 1;cactus_sprite[2][25][41] = 1;cactus_sprite[2][25][42] = 1;cactus_sprite[2][25][43] = 1;cactus_sprite[2][25][44] = 1;cactus_sprite[2][25][45] = 1;cactus_sprite[2][25][46] = 1;cactus_sprite[2][25][47] = 1;cactus_sprite[2][25][48] = 1;cactus_sprite[2][25][49] = 1;cactus_sprite[2][25][50] = 1;cactus_sprite[2][25][51] = 1;cactus_sprite[2][25][52] = 1;cactus_sprite[2][25][53] = 1;cactus_sprite[2][25][54] = 1;cactus_sprite[2][25][55] = 1;cactus_sprite[2][25][56] = 1;cactus_sprite[2][25][57] = 1;cactus_sprite[2][25][58] = 1;cactus_sprite[2][25][59] = 1;cactus_sprite[2][25][60] = 1;cactus_sprite[2][25][61] = 1;cactus_sprite[2][25][62] = 1;cactus_sprite[2][25][63] = 1;cactus_sprite[2][25][64] = 1;cactus_sprite[2][25][65] = 1;cactus_sprite[2][25][66] = 1;cactus_sprite[2][25][67] = 1;cactus_sprite[2][25][68] = 1;cactus_sprite[2][25][69] = 1;cactus_sprite[2][25][70] = 1;cactus_sprite[2][25][71] = 1;cactus_sprite[2][25][72] = 1;cactus_sprite[2][25][73] = 1;cactus_sprite[2][25][74] = 1;cactus_sprite[2][25][75] = 1;cactus_sprite[2][25][76] = 1;cactus_sprite[2][25][77] = 1;cactus_sprite[2][25][78] = 1;cactus_sprite[2][25][79] = 1;cactus_sprite[2][25][80] = 1;cactus_sprite[2][25][81] = 1;cactus_sprite[2][25][82] = 1;cactus_sprite[2][25][83] = 1;cactus_sprite[2][25][84] = 1;cactus_sprite[2][25][85] = 1;cactus_sprite[2][25][86] = 1;cactus_sprite[2][25][87] = 1;cactus_sprite[2][25][88] = 1;cactus_sprite[2][25][89] = 1;cactus_sprite[2][25][90] = 1;cactus_sprite[2][25][91] = 1;cactus_sprite[2][25][92] = 1;cactus_sprite[2][25][93] = 1;cactus_sprite[2][25][94] = 1;cactus_sprite[2][25][95] = 1;cactus_sprite[2][25][96] = 1;cactus_sprite[2][25][97] = 1;cactus_sprite[2][25][98] = 1;cactus_sprite[2][25][99] = 1;cactus_sprite[2][26][8] = 1;cactus_sprite[2][26][9] = 1;cactus_sprite[2][26][10] = 1;cactus_sprite[2][26][11] = 1;cactus_sprite[2][26][12] = 1;cactus_sprite[2][26][13] = 1;cactus_sprite[2][26][14] = 1;cactus_sprite[2][26][15] = 1;cactus_sprite[2][26][16] = 1;cactus_sprite[2][26][17] = 1;cactus_sprite[2][26][18] = 1;cactus_sprite[2][26][19] = 1;cactus_sprite[2][26][20] = 1;cactus_sprite[2][26][21] = 1;cactus_sprite[2][26][22] = 1;cactus_sprite[2][26][23] = 1;cactus_sprite[2][26][24] = 1;cactus_sprite[2][26][25] = 1;cactus_sprite[2][26][26] = 1;cactus_sprite[2][26][27] = 1;cactus_sprite[2][26][28] = 1;cactus_sprite[2][26][29] = 1;cactus_sprite[2][26][30] = 1;cactus_sprite[2][26][31] = 1;cactus_sprite[2][26][32] = 1;cactus_sprite[2][26][33] = 1;cactus_sprite[2][26][34] = 1;cactus_sprite[2][26][35] = 1;cactus_sprite[2][26][36] = 1;cactus_sprite[2][26][37] = 1;cactus_sprite[2][26][38] = 1;cactus_sprite[2][26][39] = 1;cactus_sprite[2][26][40] = 1;cactus_sprite[2][26][41] = 1;cactus_sprite[2][26][42] = 1;cactus_sprite[2][26][43] = 1;cactus_sprite[2][26][44] = 1;cactus_sprite[2][26][45] = 1;cactus_sprite[2][26][46] = 1;cactus_sprite[2][26][47] = 1;cactus_sprite[2][26][48] = 1;cactus_sprite[2][26][49] = 1;cactus_sprite[2][26][50] = 1;cactus_sprite[2][26][51] = 1;cactus_sprite[2][26][52] = 1;cactus_sprite[2][26][53] = 1;cactus_sprite[2][26][54] = 1;cactus_sprite[2][26][55] = 1;cactus_sprite[2][26][56] = 1;cactus_sprite[2][26][57] = 1;cactus_sprite[2][26][58] = 1;cactus_sprite[2][26][59] = 1;cactus_sprite[2][26][60] = 1;cactus_sprite[2][26][61] = 1;cactus_sprite[2][26][62] = 1;cactus_sprite[2][26][63] = 1;cactus_sprite[2][26][64] = 1;cactus_sprite[2][26][65] = 1;cactus_sprite[2][26][66] = 1;cactus_sprite[2][26][67] = 1;cactus_sprite[2][26][68] = 1;cactus_sprite[2][26][69] = 1;cactus_sprite[2][26][70] = 1;cactus_sprite[2][26][71] = 1;cactus_sprite[2][26][72] = 1;cactus_sprite[2][26][73] = 1;cactus_sprite[2][26][74] = 1;cactus_sprite[2][26][75] = 1;cactus_sprite[2][26][76] = 1;cactus_sprite[2][26][77] = 1;cactus_sprite[2][26][78] = 1;cactus_sprite[2][26][79] = 1;cactus_sprite[2][26][80] = 1;cactus_sprite[2][26][81] = 1;cactus_sprite[2][26][82] = 1;cactus_sprite[2][26][83] = 1;cactus_sprite[2][26][84] = 1;cactus_sprite[2][26][85] = 1;cactus_sprite[2][26][86] = 1;cactus_sprite[2][26][87] = 1;cactus_sprite[2][26][88] = 1;cactus_sprite[2][26][89] = 1;cactus_sprite[2][26][90] = 1;cactus_sprite[2][26][91] = 1;cactus_sprite[2][26][92] = 1;cactus_sprite[2][26][93] = 1;cactus_sprite[2][26][94] = 1;cactus_sprite[2][26][95] = 1;cactus_sprite[2][26][96] = 1;cactus_sprite[2][26][97] = 1;cactus_sprite[2][26][98] = 1;cactus_sprite[2][26][99] = 1;cactus_sprite[2][27][8] = 1;cactus_sprite[2][27][9] = 1;cactus_sprite[2][27][10] = 1;cactus_sprite[2][27][11] = 1;cactus_sprite[2][27][12] = 1;cactus_sprite[2][27][13] = 1;cactus_sprite[2][27][14] = 1;cactus_sprite[2][27][15] = 1;cactus_sprite[2][27][16] = 1;cactus_sprite[2][27][17] = 1;cactus_sprite[2][27][18] = 1;cactus_sprite[2][27][19] = 1;cactus_sprite[2][27][20] = 1;cactus_sprite[2][27][21] = 1;cactus_sprite[2][27][22] = 1;cactus_sprite[2][27][23] = 1;cactus_sprite[2][27][24] = 1;cactus_sprite[2][27][25] = 1;cactus_sprite[2][27][26] = 1;cactus_sprite[2][27][27] = 1;cactus_sprite[2][27][28] = 1;cactus_sprite[2][27][29] = 1;cactus_sprite[2][27][30] = 1;cactus_sprite[2][27][31] = 1;cactus_sprite[2][27][32] = 1;cactus_sprite[2][27][33] = 1;cactus_sprite[2][27][34] = 1;cactus_sprite[2][27][35] = 1;cactus_sprite[2][27][36] = 1;cactus_sprite[2][27][37] = 1;cactus_sprite[2][27][38] = 1;cactus_sprite[2][27][39] = 1;cactus_sprite[2][27][40] = 1;cactus_sprite[2][27][41] = 1;cactus_sprite[2][27][42] = 1;cactus_sprite[2][27][43] = 1;cactus_sprite[2][27][44] = 1;cactus_sprite[2][27][45] = 1;cactus_sprite[2][27][46] = 1;cactus_sprite[2][27][47] = 1;cactus_sprite[2][27][48] = 1;cactus_sprite[2][27][49] = 1;cactus_sprite[2][27][50] = 1;cactus_sprite[2][27][51] = 1;cactus_sprite[2][27][52] = 1;cactus_sprite[2][27][53] = 1;cactus_sprite[2][27][54] = 1;cactus_sprite[2][27][55] = 1;cactus_sprite[2][27][56] = 1;cactus_sprite[2][27][57] = 1;cactus_sprite[2][27][58] = 1;cactus_sprite[2][27][59] = 1;cactus_sprite[2][27][60] = 1;cactus_sprite[2][27][61] = 1;cactus_sprite[2][27][62] = 1;cactus_sprite[2][27][63] = 1;cactus_sprite[2][27][64] = 1;cactus_sprite[2][27][65] = 1;cactus_sprite[2][27][66] = 1;cactus_sprite[2][27][67] = 1;cactus_sprite[2][27][68] = 1;cactus_sprite[2][27][69] = 1;cactus_sprite[2][27][70] = 1;cactus_sprite[2][27][71] = 1;cactus_sprite[2][27][72] = 1;cactus_sprite[2][27][73] = 1;cactus_sprite[2][27][74] = 1;cactus_sprite[2][27][75] = 1;cactus_sprite[2][27][76] = 1;cactus_sprite[2][27][77] = 1;cactus_sprite[2][27][78] = 1;cactus_sprite[2][27][79] = 1;cactus_sprite[2][27][80] = 1;cactus_sprite[2][27][81] = 1;cactus_sprite[2][27][82] = 1;cactus_sprite[2][27][83] = 1;cactus_sprite[2][27][84] = 1;cactus_sprite[2][27][85] = 1;cactus_sprite[2][27][86] = 1;cactus_sprite[2][27][87] = 1;cactus_sprite[2][27][88] = 1;cactus_sprite[2][27][89] = 1;cactus_sprite[2][27][90] = 1;cactus_sprite[2][27][91] = 1;cactus_sprite[2][27][92] = 1;cactus_sprite[2][27][93] = 1;cactus_sprite[2][27][94] = 1;cactus_sprite[2][27][95] = 1;cactus_sprite[2][27][96] = 1;cactus_sprite[2][27][97] = 1;cactus_sprite[2][27][98] = 1;cactus_sprite[2][27][99] = 1;cactus_sprite[2][28][8] = 1;cactus_sprite[2][28][9] = 1;cactus_sprite[2][28][10] = 1;cactus_sprite[2][28][11] = 1;cactus_sprite[2][28][12] = 1;cactus_sprite[2][28][13] = 1;cactus_sprite[2][28][14] = 1;cactus_sprite[2][28][15] = 1;cactus_sprite[2][28][16] = 1;cactus_sprite[2][28][17] = 1;cactus_sprite[2][28][18] = 1;cactus_sprite[2][28][19] = 1;cactus_sprite[2][28][20] = 1;cactus_sprite[2][28][21] = 1;cactus_sprite[2][28][22] = 1;cactus_sprite[2][28][23] = 1;cactus_sprite[2][28][24] = 1;cactus_sprite[2][28][25] = 1;cactus_sprite[2][28][26] = 1;cactus_sprite[2][28][27] = 1;cactus_sprite[2][28][28] = 1;cactus_sprite[2][28][29] = 1;cactus_sprite[2][28][30] = 1;cactus_sprite[2][28][31] = 1;cactus_sprite[2][28][32] = 1;cactus_sprite[2][28][33] = 1;cactus_sprite[2][28][34] = 1;cactus_sprite[2][28][35] = 1;cactus_sprite[2][28][36] = 1;cactus_sprite[2][28][37] = 1;cactus_sprite[2][28][38] = 1;cactus_sprite[2][28][39] = 1;cactus_sprite[2][28][40] = 1;cactus_sprite[2][28][41] = 1;cactus_sprite[2][28][42] = 1;cactus_sprite[2][28][43] = 1;cactus_sprite[2][28][44] = 1;cactus_sprite[2][28][45] = 1;cactus_sprite[2][28][46] = 1;cactus_sprite[2][28][47] = 1;cactus_sprite[2][28][48] = 1;cactus_sprite[2][28][49] = 1;cactus_sprite[2][28][50] = 1;cactus_sprite[2][28][51] = 1;cactus_sprite[2][28][52] = 1;cactus_sprite[2][28][53] = 1;cactus_sprite[2][28][54] = 1;cactus_sprite[2][28][55] = 1;cactus_sprite[2][28][56] = 1;cactus_sprite[2][28][57] = 1;cactus_sprite[2][28][58] = 1;cactus_sprite[2][28][59] = 1;cactus_sprite[2][28][60] = 1;cactus_sprite[2][28][61] = 1;cactus_sprite[2][28][62] = 1;cactus_sprite[2][28][63] = 1;cactus_sprite[2][28][64] = 1;cactus_sprite[2][28][65] = 1;cactus_sprite[2][28][66] = 1;cactus_sprite[2][28][67] = 1;cactus_sprite[2][28][68] = 1;cactus_sprite[2][28][69] = 1;cactus_sprite[2][28][70] = 1;cactus_sprite[2][28][71] = 1;cactus_sprite[2][28][72] = 1;cactus_sprite[2][28][73] = 1;cactus_sprite[2][28][74] = 1;cactus_sprite[2][28][75] = 1;cactus_sprite[2][28][76] = 1;cactus_sprite[2][28][77] = 1;cactus_sprite[2][28][78] = 1;cactus_sprite[2][28][79] = 1;cactus_sprite[2][28][80] = 1;cactus_sprite[2][28][81] = 1;cactus_sprite[2][28][82] = 1;cactus_sprite[2][28][83] = 1;cactus_sprite[2][28][84] = 1;cactus_sprite[2][28][85] = 1;cactus_sprite[2][28][86] = 1;cactus_sprite[2][28][87] = 1;cactus_sprite[2][28][88] = 1;cactus_sprite[2][28][89] = 1;cactus_sprite[2][28][90] = 1;cactus_sprite[2][28][91] = 1;cactus_sprite[2][28][92] = 1;cactus_sprite[2][28][93] = 1;cactus_sprite[2][28][94] = 1;cactus_sprite[2][28][95] = 1;cactus_sprite[2][28][96] = 1;cactus_sprite[2][28][97] = 1;cactus_sprite[2][28][98] = 1;cactus_sprite[2][28][99] = 1;cactus_sprite[2][29][8] = 1;cactus_sprite[2][29][9] = 1;cactus_sprite[2][29][10] = 1;cactus_sprite[2][29][11] = 1;cactus_sprite[2][29][12] = 1;cactus_sprite[2][29][13] = 1;cactus_sprite[2][29][14] = 1;cactus_sprite[2][29][15] = 1;cactus_sprite[2][29][16] = 1;cactus_sprite[2][29][17] = 1;cactus_sprite[2][29][18] = 1;cactus_sprite[2][29][19] = 1;cactus_sprite[2][29][20] = 1;cactus_sprite[2][29][21] = 1;cactus_sprite[2][29][22] = 1;cactus_sprite[2][29][23] = 1;cactus_sprite[2][29][24] = 1;cactus_sprite[2][29][25] = 1;cactus_sprite[2][29][26] = 1;cactus_sprite[2][29][27] = 1;cactus_sprite[2][29][28] = 1;cactus_sprite[2][29][29] = 1;cactus_sprite[2][29][30] = 1;cactus_sprite[2][29][31] = 1;cactus_sprite[2][29][32] = 1;cactus_sprite[2][29][33] = 1;cactus_sprite[2][29][34] = 1;cactus_sprite[2][29][35] = 1;cactus_sprite[2][29][36] = 1;cactus_sprite[2][29][37] = 1;cactus_sprite[2][29][38] = 1;cactus_sprite[2][29][39] = 1;cactus_sprite[2][29][40] = 1;cactus_sprite[2][29][41] = 1;cactus_sprite[2][29][42] = 1;cactus_sprite[2][29][43] = 1;cactus_sprite[2][29][44] = 1;cactus_sprite[2][29][45] = 1;cactus_sprite[2][29][46] = 1;cactus_sprite[2][29][47] = 1;cactus_sprite[2][29][48] = 1;cactus_sprite[2][29][49] = 1;cactus_sprite[2][29][50] = 1;cactus_sprite[2][29][51] = 1;cactus_sprite[2][29][52] = 1;cactus_sprite[2][29][53] = 1;cactus_sprite[2][29][54] = 1;cactus_sprite[2][29][55] = 1;cactus_sprite[2][29][56] = 1;cactus_sprite[2][29][57] = 1;cactus_sprite[2][29][58] = 1;cactus_sprite[2][29][59] = 1;cactus_sprite[2][29][60] = 1;cactus_sprite[2][29][61] = 1;cactus_sprite[2][29][62] = 1;cactus_sprite[2][29][63] = 1;cactus_sprite[2][29][64] = 1;cactus_sprite[2][29][65] = 1;cactus_sprite[2][29][66] = 1;cactus_sprite[2][29][67] = 1;cactus_sprite[2][29][68] = 1;cactus_sprite[2][29][69] = 1;cactus_sprite[2][29][70] = 1;cactus_sprite[2][29][71] = 1;cactus_sprite[2][29][72] = 1;cactus_sprite[2][29][73] = 1;cactus_sprite[2][29][74] = 1;cactus_sprite[2][29][75] = 1;cactus_sprite[2][29][76] = 1;cactus_sprite[2][29][77] = 1;cactus_sprite[2][29][78] = 1;cactus_sprite[2][29][79] = 1;cactus_sprite[2][29][80] = 1;cactus_sprite[2][29][81] = 1;cactus_sprite[2][29][82] = 1;cactus_sprite[2][29][83] = 1;cactus_sprite[2][29][84] = 1;cactus_sprite[2][29][85] = 1;cactus_sprite[2][29][86] = 1;cactus_sprite[2][29][87] = 1;cactus_sprite[2][29][88] = 1;cactus_sprite[2][29][89] = 1;cactus_sprite[2][29][90] = 1;cactus_sprite[2][29][91] = 1;cactus_sprite[2][29][92] = 1;cactus_sprite[2][29][93] = 1;cactus_sprite[2][29][94] = 1;cactus_sprite[2][29][95] = 1;cactus_sprite[2][29][96] = 1;cactus_sprite[2][29][97] = 1;cactus_sprite[2][29][98] = 1;cactus_sprite[2][29][99] = 1;cactus_sprite[2][30][10] = 1;cactus_sprite[2][30][11] = 1;cactus_sprite[2][30][12] = 1;cactus_sprite[2][30][13] = 1;cactus_sprite[2][30][14] = 1;cactus_sprite[2][30][15] = 1;cactus_sprite[2][30][16] = 1;cactus_sprite[2][30][17] = 1;cactus_sprite[2][30][18] = 1;cactus_sprite[2][30][19] = 1;cactus_sprite[2][30][20] = 1;cactus_sprite[2][30][21] = 1;cactus_sprite[2][30][22] = 1;cactus_sprite[2][30][23] = 1;cactus_sprite[2][30][24] = 1;cactus_sprite[2][30][25] = 1;cactus_sprite[2][30][26] = 1;cactus_sprite[2][30][27] = 1;cactus_sprite[2][30][28] = 1;cactus_sprite[2][30][29] = 1;cactus_sprite[2][30][30] = 1;cactus_sprite[2][30][31] = 1;cactus_sprite[2][30][32] = 1;cactus_sprite[2][30][33] = 1;cactus_sprite[2][30][34] = 1;cactus_sprite[2][30][35] = 1;cactus_sprite[2][30][36] = 1;cactus_sprite[2][30][37] = 1;cactus_sprite[2][30][38] = 1;cactus_sprite[2][30][39] = 1;cactus_sprite[2][30][40] = 1;cactus_sprite[2][30][41] = 1;cactus_sprite[2][30][42] = 1;cactus_sprite[2][30][43] = 1;cactus_sprite[2][30][44] = 1;cactus_sprite[2][30][45] = 1;cactus_sprite[2][30][46] = 1;cactus_sprite[2][30][47] = 1;cactus_sprite[2][30][48] = 1;cactus_sprite[2][30][49] = 1;cactus_sprite[2][30][50] = 1;cactus_sprite[2][30][51] = 1;cactus_sprite[2][30][52] = 1;cactus_sprite[2][30][53] = 1;cactus_sprite[2][30][54] = 1;cactus_sprite[2][30][55] = 1;cactus_sprite[2][30][56] = 1;cactus_sprite[2][30][57] = 1;cactus_sprite[2][30][58] = 1;cactus_sprite[2][30][59] = 1;cactus_sprite[2][30][60] = 1;cactus_sprite[2][30][61] = 1;cactus_sprite[2][30][62] = 1;cactus_sprite[2][30][63] = 1;cactus_sprite[2][30][64] = 1;cactus_sprite[2][30][65] = 1;cactus_sprite[2][30][66] = 1;cactus_sprite[2][30][67] = 1;cactus_sprite[2][30][68] = 1;cactus_sprite[2][30][69] = 1;cactus_sprite[2][30][70] = 1;cactus_sprite[2][30][71] = 1;cactus_sprite[2][30][72] = 1;cactus_sprite[2][30][73] = 1;cactus_sprite[2][30][74] = 1;cactus_sprite[2][30][75] = 1;cactus_sprite[2][30][76] = 1;cactus_sprite[2][30][77] = 1;cactus_sprite[2][30][78] = 1;cactus_sprite[2][30][79] = 1;cactus_sprite[2][30][80] = 1;cactus_sprite[2][30][81] = 1;cactus_sprite[2][30][82] = 1;cactus_sprite[2][30][83] = 1;cactus_sprite[2][30][84] = 1;cactus_sprite[2][30][85] = 1;cactus_sprite[2][30][86] = 1;cactus_sprite[2][30][87] = 1;cactus_sprite[2][30][88] = 1;cactus_sprite[2][30][89] = 1;cactus_sprite[2][30][90] = 1;cactus_sprite[2][30][91] = 1;cactus_sprite[2][30][92] = 1;cactus_sprite[2][30][93] = 1;cactus_sprite[2][30][94] = 1;cactus_sprite[2][30][95] = 1;cactus_sprite[2][30][96] = 1;cactus_sprite[2][30][97] = 1;cactus_sprite[2][30][98] = 1;cactus_sprite[2][30][99] = 1;cactus_sprite[2][31][10] = 1;cactus_sprite[2][31][11] = 1;cactus_sprite[2][31][12] = 1;cactus_sprite[2][31][13] = 1;cactus_sprite[2][31][14] = 1;cactus_sprite[2][31][15] = 1;cactus_sprite[2][31][16] = 1;cactus_sprite[2][31][17] = 1;cactus_sprite[2][31][18] = 1;cactus_sprite[2][31][19] = 1;cactus_sprite[2][31][20] = 1;cactus_sprite[2][31][21] = 1;cactus_sprite[2][31][22] = 1;cactus_sprite[2][31][23] = 1;cactus_sprite[2][31][24] = 1;cactus_sprite[2][31][25] = 1;cactus_sprite[2][31][26] = 1;cactus_sprite[2][31][27] = 1;cactus_sprite[2][31][28] = 1;cactus_sprite[2][31][29] = 1;cactus_sprite[2][31][30] = 1;cactus_sprite[2][31][31] = 1;cactus_sprite[2][31][32] = 1;cactus_sprite[2][31][33] = 1;cactus_sprite[2][31][34] = 1;cactus_sprite[2][31][35] = 1;cactus_sprite[2][31][36] = 1;cactus_sprite[2][31][37] = 1;cactus_sprite[2][31][38] = 1;cactus_sprite[2][31][39] = 1;cactus_sprite[2][31][40] = 1;cactus_sprite[2][31][41] = 1;cactus_sprite[2][31][42] = 1;cactus_sprite[2][31][43] = 1;cactus_sprite[2][31][44] = 1;cactus_sprite[2][31][45] = 1;cactus_sprite[2][31][46] = 1;cactus_sprite[2][31][47] = 1;cactus_sprite[2][31][48] = 1;cactus_sprite[2][31][49] = 1;cactus_sprite[2][31][50] = 1;cactus_sprite[2][31][51] = 1;cactus_sprite[2][31][52] = 1;cactus_sprite[2][31][53] = 1;cactus_sprite[2][31][54] = 1;cactus_sprite[2][31][55] = 1;cactus_sprite[2][31][56] = 1;cactus_sprite[2][31][57] = 1;cactus_sprite[2][31][58] = 1;cactus_sprite[2][31][59] = 1;cactus_sprite[2][31][60] = 1;cactus_sprite[2][31][61] = 1;cactus_sprite[2][31][62] = 1;cactus_sprite[2][31][63] = 1;cactus_sprite[2][31][64] = 1;cactus_sprite[2][31][65] = 1;cactus_sprite[2][31][66] = 1;cactus_sprite[2][31][67] = 1;cactus_sprite[2][31][68] = 1;cactus_sprite[2][31][69] = 1;cactus_sprite[2][31][70] = 1;cactus_sprite[2][31][71] = 1;cactus_sprite[2][31][72] = 1;cactus_sprite[2][31][73] = 1;cactus_sprite[2][31][74] = 1;cactus_sprite[2][31][75] = 1;cactus_sprite[2][31][76] = 1;cactus_sprite[2][31][77] = 1;cactus_sprite[2][31][78] = 1;cactus_sprite[2][31][79] = 1;cactus_sprite[2][31][80] = 1;cactus_sprite[2][31][81] = 1;cactus_sprite[2][31][82] = 1;cactus_sprite[2][31][83] = 1;cactus_sprite[2][31][84] = 1;cactus_sprite[2][31][85] = 1;cactus_sprite[2][31][86] = 1;cactus_sprite[2][31][87] = 1;cactus_sprite[2][31][88] = 1;cactus_sprite[2][31][89] = 1;cactus_sprite[2][31][90] = 1;cactus_sprite[2][31][91] = 1;cactus_sprite[2][31][92] = 1;cactus_sprite[2][31][93] = 1;cactus_sprite[2][31][94] = 1;cactus_sprite[2][31][95] = 1;cactus_sprite[2][31][96] = 1;cactus_sprite[2][31][97] = 1;cactus_sprite[2][31][98] = 1;cactus_sprite[2][31][99] = 1;cactus_sprite[2][32][60] = 1;cactus_sprite[2][32][61] = 1;cactus_sprite[2][32][62] = 1;cactus_sprite[2][32][63] = 1;cactus_sprite[2][32][64] = 1;cactus_sprite[2][32][65] = 1;cactus_sprite[2][33][60] = 1;cactus_sprite[2][33][61] = 1;cactus_sprite[2][33][62] = 1;cactus_sprite[2][33][63] = 1;cactus_sprite[2][33][64] = 1;cactus_sprite[2][33][65] = 1;cactus_sprite[2][34][60] = 1;cactus_sprite[2][34][61] = 1;cactus_sprite[2][34][62] = 1;cactus_sprite[2][34][63] = 1;cactus_sprite[2][34][64] = 1;cactus_sprite[2][34][65] = 1;cactus_sprite[2][35][60] = 1;cactus_sprite[2][35][61] = 1;cactus_sprite[2][35][62] = 1;cactus_sprite[2][35][63] = 1;cactus_sprite[2][35][64] = 1;cactus_sprite[2][35][65] = 1;cactus_sprite[2][36][60] = 1;cactus_sprite[2][36][61] = 1;cactus_sprite[2][36][62] = 1;cactus_sprite[2][36][63] = 1;cactus_sprite[2][36][64] = 1;cactus_sprite[2][36][65] = 1;cactus_sprite[2][37][60] = 1;cactus_sprite[2][37][61] = 1;cactus_sprite[2][37][62] = 1;cactus_sprite[2][37][63] = 1;cactus_sprite[2][37][64] = 1;cactus_sprite[2][37][65] = 1;cactus_sprite[2][38][30] = 1;cactus_sprite[2][38][31] = 1;cactus_sprite[2][38][32] = 1;cactus_sprite[2][38][33] = 1;cactus_sprite[2][38][34] = 1;cactus_sprite[2][38][35] = 1;cactus_sprite[2][38][36] = 1;cactus_sprite[2][38][37] = 1;cactus_sprite[2][38][38] = 1;cactus_sprite[2][38][39] = 1;cactus_sprite[2][38][40] = 1;cactus_sprite[2][38][41] = 1;cactus_sprite[2][38][42] = 1;cactus_sprite[2][38][43] = 1;cactus_sprite[2][38][44] = 1;cactus_sprite[2][38][45] = 1;cactus_sprite[2][38][46] = 1;cactus_sprite[2][38][47] = 1;cactus_sprite[2][38][48] = 1;cactus_sprite[2][38][49] = 1;cactus_sprite[2][38][50] = 1;cactus_sprite[2][38][51] = 1;cactus_sprite[2][38][52] = 1;cactus_sprite[2][38][53] = 1;cactus_sprite[2][38][54] = 1;cactus_sprite[2][38][55] = 1;cactus_sprite[2][38][56] = 1;cactus_sprite[2][38][57] = 1;cactus_sprite[2][38][58] = 1;cactus_sprite[2][38][59] = 1;cactus_sprite[2][38][60] = 1;cactus_sprite[2][38][61] = 1;cactus_sprite[2][38][62] = 1;cactus_sprite[2][38][63] = 1;cactus_sprite[2][38][64] = 1;cactus_sprite[2][38][65] = 1;cactus_sprite[2][39][30] = 1;cactus_sprite[2][39][31] = 1;cactus_sprite[2][39][32] = 1;cactus_sprite[2][39][33] = 1;cactus_sprite[2][39][34] = 1;cactus_sprite[2][39][35] = 1;cactus_sprite[2][39][36] = 1;cactus_sprite[2][39][37] = 1;cactus_sprite[2][39][38] = 1;cactus_sprite[2][39][39] = 1;cactus_sprite[2][39][40] = 1;cactus_sprite[2][39][41] = 1;cactus_sprite[2][39][42] = 1;cactus_sprite[2][39][43] = 1;cactus_sprite[2][39][44] = 1;cactus_sprite[2][39][45] = 1;cactus_sprite[2][39][46] = 1;cactus_sprite[2][39][47] = 1;cactus_sprite[2][39][48] = 1;cactus_sprite[2][39][49] = 1;cactus_sprite[2][39][50] = 1;cactus_sprite[2][39][51] = 1;cactus_sprite[2][39][52] = 1;cactus_sprite[2][39][53] = 1;cactus_sprite[2][39][54] = 1;cactus_sprite[2][39][55] = 1;cactus_sprite[2][39][56] = 1;cactus_sprite[2][39][57] = 1;cactus_sprite[2][39][58] = 1;cactus_sprite[2][39][59] = 1;cactus_sprite[2][39][60] = 1;cactus_sprite[2][39][61] = 1;cactus_sprite[2][39][62] = 1;cactus_sprite[2][39][63] = 1;cactus_sprite[2][39][64] = 1;cactus_sprite[2][39][65] = 1;cactus_sprite[2][40][28] = 1;cactus_sprite[2][40][29] = 1;cactus_sprite[2][40][30] = 1;cactus_sprite[2][40][31] = 1;cactus_sprite[2][40][32] = 1;cactus_sprite[2][40][33] = 1;cactus_sprite[2][40][34] = 1;cactus_sprite[2][40][35] = 1;cactus_sprite[2][40][36] = 1;cactus_sprite[2][40][37] = 1;cactus_sprite[2][40][38] = 1;cactus_sprite[2][40][39] = 1;cactus_sprite[2][40][40] = 1;cactus_sprite[2][40][41] = 1;cactus_sprite[2][40][42] = 1;cactus_sprite[2][40][43] = 1;cactus_sprite[2][40][44] = 1;cactus_sprite[2][40][45] = 1;cactus_sprite[2][40][46] = 1;cactus_sprite[2][40][47] = 1;cactus_sprite[2][40][48] = 1;cactus_sprite[2][40][49] = 1;cactus_sprite[2][40][50] = 1;cactus_sprite[2][40][51] = 1;cactus_sprite[2][40][52] = 1;cactus_sprite[2][40][53] = 1;cactus_sprite[2][40][54] = 1;cactus_sprite[2][40][55] = 1;cactus_sprite[2][40][56] = 1;cactus_sprite[2][40][57] = 1;cactus_sprite[2][40][58] = 1;cactus_sprite[2][40][59] = 1;cactus_sprite[2][40][60] = 1;cactus_sprite[2][40][61] = 1;cactus_sprite[2][40][62] = 1;cactus_sprite[2][40][63] = 1;cactus_sprite[2][41][28] = 1;cactus_sprite[2][41][29] = 1;cactus_sprite[2][41][30] = 1;cactus_sprite[2][41][31] = 1;cactus_sprite[2][41][32] = 1;cactus_sprite[2][41][33] = 1;cactus_sprite[2][41][34] = 1;cactus_sprite[2][41][35] = 1;cactus_sprite[2][41][36] = 1;cactus_sprite[2][41][37] = 1;cactus_sprite[2][41][38] = 1;cactus_sprite[2][41][39] = 1;cactus_sprite[2][41][40] = 1;cactus_sprite[2][41][41] = 1;cactus_sprite[2][41][42] = 1;cactus_sprite[2][41][43] = 1;cactus_sprite[2][41][44] = 1;cactus_sprite[2][41][45] = 1;cactus_sprite[2][41][46] = 1;cactus_sprite[2][41][47] = 1;cactus_sprite[2][41][48] = 1;cactus_sprite[2][41][49] = 1;cactus_sprite[2][41][50] = 1;cactus_sprite[2][41][51] = 1;cactus_sprite[2][41][52] = 1;cactus_sprite[2][41][53] = 1;cactus_sprite[2][41][54] = 1;cactus_sprite[2][41][55] = 1;cactus_sprite[2][41][56] = 1;cactus_sprite[2][41][57] = 1;cactus_sprite[2][41][58] = 1;cactus_sprite[2][41][59] = 1;cactus_sprite[2][41][60] = 1;cactus_sprite[2][41][61] = 1;cactus_sprite[2][41][62] = 1;cactus_sprite[2][41][63] = 1;cactus_sprite[2][42][28] = 1;cactus_sprite[2][42][29] = 1;cactus_sprite[2][42][30] = 1;cactus_sprite[2][42][31] = 1;cactus_sprite[2][42][32] = 1;cactus_sprite[2][42][33] = 1;cactus_sprite[2][42][34] = 1;cactus_sprite[2][42][35] = 1;cactus_sprite[2][42][36] = 1;cactus_sprite[2][42][37] = 1;cactus_sprite[2][42][38] = 1;cactus_sprite[2][42][39] = 1;cactus_sprite[2][42][40] = 1;cactus_sprite[2][42][41] = 1;cactus_sprite[2][42][42] = 1;cactus_sprite[2][42][43] = 1;cactus_sprite[2][42][44] = 1;cactus_sprite[2][42][45] = 1;cactus_sprite[2][42][46] = 1;cactus_sprite[2][42][47] = 1;cactus_sprite[2][42][48] = 1;cactus_sprite[2][42][49] = 1;cactus_sprite[2][42][50] = 1;cactus_sprite[2][42][51] = 1;cactus_sprite[2][42][52] = 1;cactus_sprite[2][42][53] = 1;cactus_sprite[2][42][54] = 1;cactus_sprite[2][42][55] = 1;cactus_sprite[2][42][56] = 1;cactus_sprite[2][42][57] = 1;cactus_sprite[2][42][58] = 1;cactus_sprite[2][42][59] = 1;cactus_sprite[2][42][60] = 1;cactus_sprite[2][42][61] = 1;cactus_sprite[2][43][28] = 1;cactus_sprite[2][43][29] = 1;cactus_sprite[2][43][30] = 1;cactus_sprite[2][43][31] = 1;cactus_sprite[2][43][32] = 1;cactus_sprite[2][43][33] = 1;cactus_sprite[2][43][34] = 1;cactus_sprite[2][43][35] = 1;cactus_sprite[2][43][36] = 1;cactus_sprite[2][43][37] = 1;cactus_sprite[2][43][38] = 1;cactus_sprite[2][43][39] = 1;cactus_sprite[2][43][40] = 1;cactus_sprite[2][43][41] = 1;cactus_sprite[2][43][42] = 1;cactus_sprite[2][43][43] = 1;cactus_sprite[2][43][44] = 1;cactus_sprite[2][43][45] = 1;cactus_sprite[2][43][46] = 1;cactus_sprite[2][43][47] = 1;cactus_sprite[2][43][48] = 1;cactus_sprite[2][43][49] = 1;cactus_sprite[2][43][50] = 1;cactus_sprite[2][43][51] = 1;cactus_sprite[2][43][52] = 1;cactus_sprite[2][43][53] = 1;cactus_sprite[2][43][54] = 1;cactus_sprite[2][43][55] = 1;cactus_sprite[2][43][56] = 1;cactus_sprite[2][43][57] = 1;cactus_sprite[2][43][58] = 1;cactus_sprite[2][43][59] = 1;cactus_sprite[2][43][60] = 1;cactus_sprite[2][43][61] = 1;cactus_sprite[2][44][30] = 1;cactus_sprite[2][44][31] = 1;cactus_sprite[2][44][32] = 1;cactus_sprite[2][44][33] = 1;cactus_sprite[2][44][34] = 1;cactus_sprite[2][44][35] = 1;cactus_sprite[2][44][36] = 1;cactus_sprite[2][44][37] = 1;cactus_sprite[2][44][38] = 1;cactus_sprite[2][44][39] = 1;cactus_sprite[2][44][40] = 1;cactus_sprite[2][44][41] = 1;cactus_sprite[2][44][42] = 1;cactus_sprite[2][44][43] = 1;cactus_sprite[2][44][44] = 1;cactus_sprite[2][44][45] = 1;cactus_sprite[2][44][46] = 1;cactus_sprite[2][44][47] = 1;cactus_sprite[2][44][48] = 1;cactus_sprite[2][44][49] = 1;cactus_sprite[2][44][50] = 1;cactus_sprite[2][44][51] = 1;cactus_sprite[2][44][52] = 1;cactus_sprite[2][44][53] = 1;cactus_sprite[2][44][54] = 1;cactus_sprite[2][44][55] = 1;cactus_sprite[2][44][56] = 1;cactus_sprite[2][44][57] = 1;cactus_sprite[2][44][58] = 1;cactus_sprite[2][44][59] = 1;cactus_sprite[2][45][30] = 1;cactus_sprite[2][45][31] = 1;cactus_sprite[2][45][32] = 1;cactus_sprite[2][45][33] = 1;cactus_sprite[2][45][34] = 1;cactus_sprite[2][45][35] = 1;cactus_sprite[2][45][36] = 1;cactus_sprite[2][45][37] = 1;cactus_sprite[2][45][38] = 1;cactus_sprite[2][45][39] = 1;cactus_sprite[2][45][40] = 1;cactus_sprite[2][45][41] = 1;cactus_sprite[2][45][42] = 1;cactus_sprite[2][45][43] = 1;cactus_sprite[2][45][44] = 1;cactus_sprite[2][45][45] = 1;cactus_sprite[2][45][46] = 1;cactus_sprite[2][45][47] = 1;cactus_sprite[2][45][48] = 1;cactus_sprite[2][45][49] = 1;cactus_sprite[2][45][50] = 1;cactus_sprite[2][45][51] = 1;cactus_sprite[2][45][52] = 1;cactus_sprite[2][45][53] = 1;cactus_sprite[2][45][54] = 1;cactus_sprite[2][45][55] = 1;cactus_sprite[2][45][56] = 1;cactus_sprite[2][45][57] = 1;cactus_sprite[2][45][58] = 1;cactus_sprite[2][45][59] = 1;
	cactus_sprite[3][2][32] = 1;cactus_sprite[3][2][33] = 1;cactus_sprite[3][2][34] = 1;cactus_sprite[3][2][35] = 1;cactus_sprite[3][2][36] = 1;cactus_sprite[3][2][37] = 1;cactus_sprite[3][2][38] = 1;cactus_sprite[3][2][39] = 1;cactus_sprite[3][2][40] = 1;cactus_sprite[3][2][41] = 1;cactus_sprite[3][2][42] = 1;cactus_sprite[3][2][43] = 1;cactus_sprite[3][2][44] = 1;cactus_sprite[3][2][45] = 1;cactus_sprite[3][2][46] = 1;cactus_sprite[3][2][47] = 1;cactus_sprite[3][2][48] = 1;cactus_sprite[3][2][49] = 1;cactus_sprite[3][2][50] = 1;cactus_sprite[3][2][51] = 1;cactus_sprite[3][2][52] = 1;cactus_sprite[3][2][53] = 1;cactus_sprite[3][2][54] = 1;cactus_sprite[3][2][55] = 1;cactus_sprite[3][2][56] = 1;cactus_sprite[3][2][57] = 1;cactus_sprite[3][2][58] = 1;cactus_sprite[3][2][59] = 1;cactus_sprite[3][2][60] = 1;cactus_sprite[3][2][61] = 1;cactus_sprite[3][3][32] = 1;cactus_sprite[3][3][33] = 1;cactus_sprite[3][3][34] = 1;cactus_sprite[3][3][35] = 1;cactus_sprite[3][3][36] = 1;cactus_sprite[3][3][37] = 1;cactus_sprite[3][3][38] = 1;cactus_sprite[3][3][39] = 1;cactus_sprite[3][3][40] = 1;cactus_sprite[3][3][41] = 1;cactus_sprite[3][3][42] = 1;cactus_sprite[3][3][43] = 1;cactus_sprite[3][3][44] = 1;cactus_sprite[3][3][45] = 1;cactus_sprite[3][3][46] = 1;cactus_sprite[3][3][47] = 1;cactus_sprite[3][3][48] = 1;cactus_sprite[3][3][49] = 1;cactus_sprite[3][3][50] = 1;cactus_sprite[3][3][51] = 1;cactus_sprite[3][3][52] = 1;cactus_sprite[3][3][53] = 1;cactus_sprite[3][3][54] = 1;cactus_sprite[3][3][55] = 1;cactus_sprite[3][3][56] = 1;cactus_sprite[3][3][57] = 1;cactus_sprite[3][3][58] = 1;cactus_sprite[3][3][59] = 1;cactus_sprite[3][3][60] = 1;cactus_sprite[3][3][61] = 1;cactus_sprite[3][4][30] = 1;cactus_sprite[3][4][31] = 1;cactus_sprite[3][4][32] = 1;cactus_sprite[3][4][33] = 1;cactus_sprite[3][4][34] = 1;cactus_sprite[3][4][35] = 1;cactus_sprite[3][4][36] = 1;cactus_sprite[3][4][37] = 1;cactus_sprite[3][4][38] = 1;cactus_sprite[3][4][39] = 1;cactus_sprite[3][4][40] = 1;cactus_sprite[3][4][41] = 1;cactus_sprite[3][4][42] = 1;cactus_sprite[3][4][43] = 1;cactus_sprite[3][4][44] = 1;cactus_sprite[3][4][45] = 1;cactus_sprite[3][4][46] = 1;cactus_sprite[3][4][47] = 1;cactus_sprite[3][4][48] = 1;cactus_sprite[3][4][49] = 1;cactus_sprite[3][4][50] = 1;cactus_sprite[3][4][51] = 1;cactus_sprite[3][4][52] = 1;cactus_sprite[3][4][53] = 1;cactus_sprite[3][4][54] = 1;cactus_sprite[3][4][55] = 1;cactus_sprite[3][4][56] = 1;cactus_sprite[3][4][57] = 1;cactus_sprite[3][4][58] = 1;cactus_sprite[3][4][59] = 1;cactus_sprite[3][4][60] = 1;cactus_sprite[3][4][61] = 1;cactus_sprite[3][4][62] = 1;cactus_sprite[3][4][63] = 1;cactus_sprite[3][5][30] = 1;cactus_sprite[3][5][31] = 1;cactus_sprite[3][5][32] = 1;cactus_sprite[3][5][33] = 1;cactus_sprite[3][5][34] = 1;cactus_sprite[3][5][35] = 1;cactus_sprite[3][5][36] = 1;cactus_sprite[3][5][37] = 1;cactus_sprite[3][5][38] = 1;cactus_sprite[3][5][39] = 1;cactus_sprite[3][5][40] = 1;cactus_sprite[3][5][41] = 1;cactus_sprite[3][5][42] = 1;cactus_sprite[3][5][43] = 1;cactus_sprite[3][5][44] = 1;cactus_sprite[3][5][45] = 1;cactus_sprite[3][5][46] = 1;cactus_sprite[3][5][47] = 1;cactus_sprite[3][5][48] = 1;cactus_sprite[3][5][49] = 1;cactus_sprite[3][5][50] = 1;cactus_sprite[3][5][51] = 1;cactus_sprite[3][5][52] = 1;cactus_sprite[3][5][53] = 1;cactus_sprite[3][5][54] = 1;cactus_sprite[3][5][55] = 1;cactus_sprite[3][5][56] = 1;cactus_sprite[3][5][57] = 1;cactus_sprite[3][5][58] = 1;cactus_sprite[3][5][59] = 1;cactus_sprite[3][5][60] = 1;cactus_sprite[3][5][61] = 1;cactus_sprite[3][5][62] = 1;cactus_sprite[3][5][63] = 1;cactus_sprite[3][6][30] = 1;cactus_sprite[3][6][31] = 1;cactus_sprite[3][6][32] = 1;cactus_sprite[3][6][33] = 1;cactus_sprite[3][6][34] = 1;cactus_sprite[3][6][35] = 1;cactus_sprite[3][6][36] = 1;cactus_sprite[3][6][37] = 1;cactus_sprite[3][6][38] = 1;cactus_sprite[3][6][39] = 1;cactus_sprite[3][6][40] = 1;cactus_sprite[3][6][41] = 1;cactus_sprite[3][6][42] = 1;cactus_sprite[3][6][43] = 1;cactus_sprite[3][6][44] = 1;cactus_sprite[3][6][45] = 1;cactus_sprite[3][6][46] = 1;cactus_sprite[3][6][47] = 1;cactus_sprite[3][6][48] = 1;cactus_sprite[3][6][49] = 1;cactus_sprite[3][6][50] = 1;cactus_sprite[3][6][51] = 1;cactus_sprite[3][6][52] = 1;cactus_sprite[3][6][53] = 1;cactus_sprite[3][6][54] = 1;cactus_sprite[3][6][55] = 1;cactus_sprite[3][6][56] = 1;cactus_sprite[3][6][57] = 1;cactus_sprite[3][6][58] = 1;cactus_sprite[3][6][59] = 1;cactus_sprite[3][6][60] = 1;cactus_sprite[3][6][61] = 1;cactus_sprite[3][6][62] = 1;cactus_sprite[3][6][63] = 1;cactus_sprite[3][6][64] = 1;cactus_sprite[3][6][65] = 1;cactus_sprite[3][7][30] = 1;cactus_sprite[3][7][31] = 1;cactus_sprite[3][7][32] = 1;cactus_sprite[3][7][33] = 1;cactus_sprite[3][7][34] = 1;cactus_sprite[3][7][35] = 1;cactus_sprite[3][7][36] = 1;cactus_sprite[3][7][37] = 1;cactus_sprite[3][7][38] = 1;cactus_sprite[3][7][39] = 1;cactus_sprite[3][7][40] = 1;cactus_sprite[3][7][41] = 1;cactus_sprite[3][7][42] = 1;cactus_sprite[3][7][43] = 1;cactus_sprite[3][7][44] = 1;cactus_sprite[3][7][45] = 1;cactus_sprite[3][7][46] = 1;cactus_sprite[3][7][47] = 1;cactus_sprite[3][7][48] = 1;cactus_sprite[3][7][49] = 1;cactus_sprite[3][7][50] = 1;cactus_sprite[3][7][51] = 1;cactus_sprite[3][7][52] = 1;cactus_sprite[3][7][53] = 1;cactus_sprite[3][7][54] = 1;cactus_sprite[3][7][55] = 1;cactus_sprite[3][7][56] = 1;cactus_sprite[3][7][57] = 1;cactus_sprite[3][7][58] = 1;cactus_sprite[3][7][59] = 1;cactus_sprite[3][7][60] = 1;cactus_sprite[3][7][61] = 1;cactus_sprite[3][7][62] = 1;cactus_sprite[3][7][63] = 1;cactus_sprite[3][7][64] = 1;cactus_sprite[3][7][65] = 1;cactus_sprite[3][8][30] = 1;cactus_sprite[3][8][31] = 1;cactus_sprite[3][8][32] = 1;cactus_sprite[3][8][33] = 1;cactus_sprite[3][8][34] = 1;cactus_sprite[3][8][35] = 1;cactus_sprite[3][8][36] = 1;cactus_sprite[3][8][37] = 1;cactus_sprite[3][8][38] = 1;cactus_sprite[3][8][39] = 1;cactus_sprite[3][8][40] = 1;cactus_sprite[3][8][41] = 1;cactus_sprite[3][8][42] = 1;cactus_sprite[3][8][43] = 1;cactus_sprite[3][8][44] = 1;cactus_sprite[3][8][45] = 1;cactus_sprite[3][8][46] = 1;cactus_sprite[3][8][47] = 1;cactus_sprite[3][8][48] = 1;cactus_sprite[3][8][49] = 1;cactus_sprite[3][8][50] = 1;cactus_sprite[3][8][51] = 1;cactus_sprite[3][8][52] = 1;cactus_sprite[3][8][53] = 1;cactus_sprite[3][8][54] = 1;cactus_sprite[3][8][55] = 1;cactus_sprite[3][8][56] = 1;cactus_sprite[3][8][57] = 1;cactus_sprite[3][8][58] = 1;cactus_sprite[3][8][59] = 1;cactus_sprite[3][8][60] = 1;cactus_sprite[3][8][61] = 1;cactus_sprite[3][8][62] = 1;cactus_sprite[3][8][63] = 1;cactus_sprite[3][8][64] = 1;cactus_sprite[3][8][65] = 1;cactus_sprite[3][8][66] = 1;cactus_sprite[3][8][67] = 1;cactus_sprite[3][9][30] = 1;cactus_sprite[3][9][31] = 1;cactus_sprite[3][9][32] = 1;cactus_sprite[3][9][33] = 1;cactus_sprite[3][9][34] = 1;cactus_sprite[3][9][35] = 1;cactus_sprite[3][9][36] = 1;cactus_sprite[3][9][37] = 1;cactus_sprite[3][9][38] = 1;cactus_sprite[3][9][39] = 1;cactus_sprite[3][9][40] = 1;cactus_sprite[3][9][41] = 1;cactus_sprite[3][9][42] = 1;cactus_sprite[3][9][43] = 1;cactus_sprite[3][9][44] = 1;cactus_sprite[3][9][45] = 1;cactus_sprite[3][9][46] = 1;cactus_sprite[3][9][47] = 1;cactus_sprite[3][9][48] = 1;cactus_sprite[3][9][49] = 1;cactus_sprite[3][9][50] = 1;cactus_sprite[3][9][51] = 1;cactus_sprite[3][9][52] = 1;cactus_sprite[3][9][53] = 1;cactus_sprite[3][9][54] = 1;cactus_sprite[3][9][55] = 1;cactus_sprite[3][9][56] = 1;cactus_sprite[3][9][57] = 1;cactus_sprite[3][9][58] = 1;cactus_sprite[3][9][59] = 1;cactus_sprite[3][9][60] = 1;cactus_sprite[3][9][61] = 1;cactus_sprite[3][9][62] = 1;cactus_sprite[3][9][63] = 1;cactus_sprite[3][9][64] = 1;cactus_sprite[3][9][65] = 1;cactus_sprite[3][9][66] = 1;cactus_sprite[3][9][67] = 1;cactus_sprite[3][10][32] = 1;cactus_sprite[3][10][33] = 1;cactus_sprite[3][10][34] = 1;cactus_sprite[3][10][35] = 1;cactus_sprite[3][10][36] = 1;cactus_sprite[3][10][37] = 1;cactus_sprite[3][10][38] = 1;cactus_sprite[3][10][39] = 1;cactus_sprite[3][10][40] = 1;cactus_sprite[3][10][41] = 1;cactus_sprite[3][10][42] = 1;cactus_sprite[3][10][43] = 1;cactus_sprite[3][10][44] = 1;cactus_sprite[3][10][45] = 1;cactus_sprite[3][10][46] = 1;cactus_sprite[3][10][47] = 1;cactus_sprite[3][10][48] = 1;cactus_sprite[3][10][49] = 1;cactus_sprite[3][10][50] = 1;cactus_sprite[3][10][51] = 1;cactus_sprite[3][10][52] = 1;cactus_sprite[3][10][53] = 1;cactus_sprite[3][10][54] = 1;cactus_sprite[3][10][55] = 1;cactus_sprite[3][10][56] = 1;cactus_sprite[3][10][57] = 1;cactus_sprite[3][10][58] = 1;cactus_sprite[3][10][59] = 1;cactus_sprite[3][10][60] = 1;cactus_sprite[3][10][61] = 1;cactus_sprite[3][10][62] = 1;cactus_sprite[3][10][63] = 1;cactus_sprite[3][10][64] = 1;cactus_sprite[3][10][65] = 1;cactus_sprite[3][10][66] = 1;cactus_sprite[3][10][67] = 1;cactus_sprite[3][10][68] = 1;cactus_sprite[3][10][69] = 1;cactus_sprite[3][11][32] = 1;cactus_sprite[3][11][33] = 1;cactus_sprite[3][11][34] = 1;cactus_sprite[3][11][35] = 1;cactus_sprite[3][11][36] = 1;cactus_sprite[3][11][37] = 1;cactus_sprite[3][11][38] = 1;cactus_sprite[3][11][39] = 1;cactus_sprite[3][11][40] = 1;cactus_sprite[3][11][41] = 1;cactus_sprite[3][11][42] = 1;cactus_sprite[3][11][43] = 1;cactus_sprite[3][11][44] = 1;cactus_sprite[3][11][45] = 1;cactus_sprite[3][11][46] = 1;cactus_sprite[3][11][47] = 1;cactus_sprite[3][11][48] = 1;cactus_sprite[3][11][49] = 1;cactus_sprite[3][11][50] = 1;cactus_sprite[3][11][51] = 1;cactus_sprite[3][11][52] = 1;cactus_sprite[3][11][53] = 1;cactus_sprite[3][11][54] = 1;cactus_sprite[3][11][55] = 1;cactus_sprite[3][11][56] = 1;cactus_sprite[3][11][57] = 1;cactus_sprite[3][11][58] = 1;cactus_sprite[3][11][59] = 1;cactus_sprite[3][11][60] = 1;cactus_sprite[3][11][61] = 1;cactus_sprite[3][11][62] = 1;cactus_sprite[3][11][63] = 1;cactus_sprite[3][11][64] = 1;cactus_sprite[3][11][65] = 1;cactus_sprite[3][11][66] = 1;cactus_sprite[3][11][67] = 1;cactus_sprite[3][11][68] = 1;cactus_sprite[3][11][69] = 1;cactus_sprite[3][12][60] = 1;cactus_sprite[3][12][61] = 1;cactus_sprite[3][12][62] = 1;cactus_sprite[3][12][63] = 1;cactus_sprite[3][12][64] = 1;cactus_sprite[3][12][65] = 1;cactus_sprite[3][12][66] = 1;cactus_sprite[3][12][67] = 1;cactus_sprite[3][12][68] = 1;cactus_sprite[3][12][69] = 1;cactus_sprite[3][13][60] = 1;cactus_sprite[3][13][61] = 1;cactus_sprite[3][13][62] = 1;cactus_sprite[3][13][63] = 1;cactus_sprite[3][13][64] = 1;cactus_sprite[3][13][65] = 1;cactus_sprite[3][13][66] = 1;cactus_sprite[3][13][67] = 1;cactus_sprite[3][13][68] = 1;cactus_sprite[3][13][69] = 1;cactus_sprite[3][14][60] = 1;cactus_sprite[3][14][61] = 1;cactus_sprite[3][14][62] = 1;cactus_sprite[3][14][63] = 1;cactus_sprite[3][14][64] = 1;cactus_sprite[3][14][65] = 1;cactus_sprite[3][14][66] = 1;cactus_sprite[3][14][67] = 1;cactus_sprite[3][14][68] = 1;cactus_sprite[3][14][69] = 1;cactus_sprite[3][15][60] = 1;cactus_sprite[3][15][61] = 1;cactus_sprite[3][15][62] = 1;cactus_sprite[3][15][63] = 1;cactus_sprite[3][15][64] = 1;cactus_sprite[3][15][65] = 1;cactus_sprite[3][15][66] = 1;cactus_sprite[3][15][67] = 1;cactus_sprite[3][15][68] = 1;cactus_sprite[3][15][69] = 1;cactus_sprite[3][16][60] = 1;cactus_sprite[3][16][61] = 1;cactus_sprite[3][16][62] = 1;cactus_sprite[3][16][63] = 1;cactus_sprite[3][16][64] = 1;cactus_sprite[3][16][65] = 1;cactus_sprite[3][16][66] = 1;cactus_sprite[3][16][67] = 1;cactus_sprite[3][16][68] = 1;cactus_sprite[3][16][69] = 1;cactus_sprite[3][17][60] = 1;cactus_sprite[3][17][61] = 1;cactus_sprite[3][17][62] = 1;cactus_sprite[3][17][63] = 1;cactus_sprite[3][17][64] = 1;cactus_sprite[3][17][65] = 1;cactus_sprite[3][17][66] = 1;cactus_sprite[3][17][67] = 1;cactus_sprite[3][17][68] = 1;cactus_sprite[3][17][69] = 1;cactus_sprite[3][18][8] = 1;cactus_sprite[3][18][9] = 1;cactus_sprite[3][18][10] = 1;cactus_sprite[3][18][11] = 1;cactus_sprite[3][18][12] = 1;cactus_sprite[3][18][13] = 1;cactus_sprite[3][18][14] = 1;cactus_sprite[3][18][15] = 1;cactus_sprite[3][18][16] = 1;cactus_sprite[3][18][17] = 1;cactus_sprite[3][18][18] = 1;cactus_sprite[3][18][19] = 1;cactus_sprite[3][18][20] = 1;cactus_sprite[3][18][21] = 1;cactus_sprite[3][18][22] = 1;cactus_sprite[3][18][23] = 1;cactus_sprite[3][18][24] = 1;cactus_sprite[3][18][25] = 1;cactus_sprite[3][18][26] = 1;cactus_sprite[3][18][27] = 1;cactus_sprite[3][18][28] = 1;cactus_sprite[3][18][29] = 1;cactus_sprite[3][18][30] = 1;cactus_sprite[3][18][31] = 1;cactus_sprite[3][18][32] = 1;cactus_sprite[3][18][33] = 1;cactus_sprite[3][18][34] = 1;cactus_sprite[3][18][35] = 1;cactus_sprite[3][18][36] = 1;cactus_sprite[3][18][37] = 1;cactus_sprite[3][18][38] = 1;cactus_sprite[3][18][39] = 1;cactus_sprite[3][18][40] = 1;cactus_sprite[3][18][41] = 1;cactus_sprite[3][18][42] = 1;cactus_sprite[3][18][43] = 1;cactus_sprite[3][18][44] = 1;cactus_sprite[3][18][45] = 1;cactus_sprite[3][18][46] = 1;cactus_sprite[3][18][47] = 1;cactus_sprite[3][18][48] = 1;cactus_sprite[3][18][49] = 1;cactus_sprite[3][18][50] = 1;cactus_sprite[3][18][51] = 1;cactus_sprite[3][18][52] = 1;cactus_sprite[3][18][53] = 1;cactus_sprite[3][18][54] = 1;cactus_sprite[3][18][55] = 1;cactus_sprite[3][18][56] = 1;cactus_sprite[3][18][57] = 1;cactus_sprite[3][18][58] = 1;cactus_sprite[3][18][59] = 1;cactus_sprite[3][18][60] = 1;cactus_sprite[3][18][61] = 1;cactus_sprite[3][18][62] = 1;cactus_sprite[3][18][63] = 1;cactus_sprite[3][18][64] = 1;cactus_sprite[3][18][65] = 1;cactus_sprite[3][18][66] = 1;cactus_sprite[3][18][67] = 1;cactus_sprite[3][18][68] = 1;cactus_sprite[3][18][69] = 1;cactus_sprite[3][18][70] = 1;cactus_sprite[3][18][71] = 1;cactus_sprite[3][18][72] = 1;cactus_sprite[3][18][73] = 1;cactus_sprite[3][18][74] = 1;cactus_sprite[3][18][75] = 1;cactus_sprite[3][18][76] = 1;cactus_sprite[3][18][77] = 1;cactus_sprite[3][18][78] = 1;cactus_sprite[3][18][79] = 1;cactus_sprite[3][18][80] = 1;cactus_sprite[3][18][81] = 1;cactus_sprite[3][18][82] = 1;cactus_sprite[3][18][83] = 1;cactus_sprite[3][18][84] = 1;cactus_sprite[3][18][85] = 1;cactus_sprite[3][18][86] = 1;cactus_sprite[3][18][87] = 1;cactus_sprite[3][18][88] = 1;cactus_sprite[3][18][89] = 1;cactus_sprite[3][18][90] = 1;cactus_sprite[3][18][91] = 1;cactus_sprite[3][18][92] = 1;cactus_sprite[3][18][93] = 1;cactus_sprite[3][18][94] = 1;cactus_sprite[3][18][95] = 1;cactus_sprite[3][18][96] = 1;cactus_sprite[3][18][97] = 1;cactus_sprite[3][18][98] = 1;cactus_sprite[3][18][99] = 1;cactus_sprite[3][19][8] = 1;cactus_sprite[3][19][9] = 1;cactus_sprite[3][19][10] = 1;cactus_sprite[3][19][11] = 1;cactus_sprite[3][19][12] = 1;cactus_sprite[3][19][13] = 1;cactus_sprite[3][19][14] = 1;cactus_sprite[3][19][15] = 1;cactus_sprite[3][19][16] = 1;cactus_sprite[3][19][17] = 1;cactus_sprite[3][19][18] = 1;cactus_sprite[3][19][19] = 1;cactus_sprite[3][19][20] = 1;cactus_sprite[3][19][21] = 1;cactus_sprite[3][19][22] = 1;cactus_sprite[3][19][23] = 1;cactus_sprite[3][19][24] = 1;cactus_sprite[3][19][25] = 1;cactus_sprite[3][19][26] = 1;cactus_sprite[3][19][27] = 1;cactus_sprite[3][19][28] = 1;cactus_sprite[3][19][29] = 1;cactus_sprite[3][19][30] = 1;cactus_sprite[3][19][31] = 1;cactus_sprite[3][19][32] = 1;cactus_sprite[3][19][33] = 1;cactus_sprite[3][19][34] = 1;cactus_sprite[3][19][35] = 1;cactus_sprite[3][19][36] = 1;cactus_sprite[3][19][37] = 1;cactus_sprite[3][19][38] = 1;cactus_sprite[3][19][39] = 1;cactus_sprite[3][19][40] = 1;cactus_sprite[3][19][41] = 1;cactus_sprite[3][19][42] = 1;cactus_sprite[3][19][43] = 1;cactus_sprite[3][19][44] = 1;cactus_sprite[3][19][45] = 1;cactus_sprite[3][19][46] = 1;cactus_sprite[3][19][47] = 1;cactus_sprite[3][19][48] = 1;cactus_sprite[3][19][49] = 1;cactus_sprite[3][19][50] = 1;cactus_sprite[3][19][51] = 1;cactus_sprite[3][19][52] = 1;cactus_sprite[3][19][53] = 1;cactus_sprite[3][19][54] = 1;cactus_sprite[3][19][55] = 1;cactus_sprite[3][19][56] = 1;cactus_sprite[3][19][57] = 1;cactus_sprite[3][19][58] = 1;cactus_sprite[3][19][59] = 1;cactus_sprite[3][19][60] = 1;cactus_sprite[3][19][61] = 1;cactus_sprite[3][19][62] = 1;cactus_sprite[3][19][63] = 1;cactus_sprite[3][19][64] = 1;cactus_sprite[3][19][65] = 1;cactus_sprite[3][19][66] = 1;cactus_sprite[3][19][67] = 1;cactus_sprite[3][19][68] = 1;cactus_sprite[3][19][69] = 1;cactus_sprite[3][19][70] = 1;cactus_sprite[3][19][71] = 1;cactus_sprite[3][19][72] = 1;cactus_sprite[3][19][73] = 1;cactus_sprite[3][19][74] = 1;cactus_sprite[3][19][75] = 1;cactus_sprite[3][19][76] = 1;cactus_sprite[3][19][77] = 1;cactus_sprite[3][19][78] = 1;cactus_sprite[3][19][79] = 1;cactus_sprite[3][19][80] = 1;cactus_sprite[3][19][81] = 1;cactus_sprite[3][19][82] = 1;cactus_sprite[3][19][83] = 1;cactus_sprite[3][19][84] = 1;cactus_sprite[3][19][85] = 1;cactus_sprite[3][19][86] = 1;cactus_sprite[3][19][87] = 1;cactus_sprite[3][19][88] = 1;cactus_sprite[3][19][89] = 1;cactus_sprite[3][19][90] = 1;cactus_sprite[3][19][91] = 1;cactus_sprite[3][19][92] = 1;cactus_sprite[3][19][93] = 1;cactus_sprite[3][19][94] = 1;cactus_sprite[3][19][95] = 1;cactus_sprite[3][19][96] = 1;cactus_sprite[3][19][97] = 1;cactus_sprite[3][19][98] = 1;cactus_sprite[3][19][99] = 1;cactus_sprite[3][20][6] = 1;cactus_sprite[3][20][7] = 1;cactus_sprite[3][20][8] = 1;cactus_sprite[3][20][9] = 1;cactus_sprite[3][20][10] = 1;cactus_sprite[3][20][11] = 1;cactus_sprite[3][20][12] = 1;cactus_sprite[3][20][13] = 1;cactus_sprite[3][20][14] = 1;cactus_sprite[3][20][15] = 1;cactus_sprite[3][20][16] = 1;cactus_sprite[3][20][17] = 1;cactus_sprite[3][20][18] = 1;cactus_sprite[3][20][19] = 1;cactus_sprite[3][20][20] = 1;cactus_sprite[3][20][21] = 1;cactus_sprite[3][20][22] = 1;cactus_sprite[3][20][23] = 1;cactus_sprite[3][20][24] = 1;cactus_sprite[3][20][25] = 1;cactus_sprite[3][20][26] = 1;cactus_sprite[3][20][27] = 1;cactus_sprite[3][20][28] = 1;cactus_sprite[3][20][29] = 1;cactus_sprite[3][20][30] = 1;cactus_sprite[3][20][31] = 1;cactus_sprite[3][20][32] = 1;cactus_sprite[3][20][33] = 1;cactus_sprite[3][20][34] = 1;cactus_sprite[3][20][35] = 1;cactus_sprite[3][20][36] = 1;cactus_sprite[3][20][37] = 1;cactus_sprite[3][20][38] = 1;cactus_sprite[3][20][39] = 1;cactus_sprite[3][20][40] = 1;cactus_sprite[3][20][41] = 1;cactus_sprite[3][20][42] = 1;cactus_sprite[3][20][43] = 1;cactus_sprite[3][20][44] = 1;cactus_sprite[3][20][45] = 1;cactus_sprite[3][20][46] = 1;cactus_sprite[3][20][47] = 1;cactus_sprite[3][20][48] = 1;cactus_sprite[3][20][49] = 1;cactus_sprite[3][20][50] = 1;cactus_sprite[3][20][51] = 1;cactus_sprite[3][20][52] = 1;cactus_sprite[3][20][53] = 1;cactus_sprite[3][20][54] = 1;cactus_sprite[3][20][55] = 1;cactus_sprite[3][20][56] = 1;cactus_sprite[3][20][57] = 1;cactus_sprite[3][20][58] = 1;cactus_sprite[3][20][59] = 1;cactus_sprite[3][20][60] = 1;cactus_sprite[3][20][61] = 1;cactus_sprite[3][20][62] = 1;cactus_sprite[3][20][63] = 1;cactus_sprite[3][20][64] = 1;cactus_sprite[3][20][65] = 1;cactus_sprite[3][20][66] = 1;cactus_sprite[3][20][67] = 1;cactus_sprite[3][20][68] = 1;cactus_sprite[3][20][69] = 1;cactus_sprite[3][20][70] = 1;cactus_sprite[3][20][71] = 1;cactus_sprite[3][20][72] = 1;cactus_sprite[3][20][73] = 1;cactus_sprite[3][20][74] = 1;cactus_sprite[3][20][75] = 1;cactus_sprite[3][20][76] = 1;cactus_sprite[3][20][77] = 1;cactus_sprite[3][20][78] = 1;cactus_sprite[3][20][79] = 1;cactus_sprite[3][20][80] = 1;cactus_sprite[3][20][81] = 1;cactus_sprite[3][20][82] = 1;cactus_sprite[3][20][83] = 1;cactus_sprite[3][20][84] = 1;cactus_sprite[3][20][85] = 1;cactus_sprite[3][20][86] = 1;cactus_sprite[3][20][87] = 1;cactus_sprite[3][20][88] = 1;cactus_sprite[3][20][89] = 1;cactus_sprite[3][20][90] = 1;cactus_sprite[3][20][91] = 1;cactus_sprite[3][20][92] = 1;cactus_sprite[3][20][93] = 1;cactus_sprite[3][20][94] = 1;cactus_sprite[3][20][95] = 1;cactus_sprite[3][20][96] = 1;cactus_sprite[3][20][97] = 1;cactus_sprite[3][20][98] = 1;cactus_sprite[3][20][99] = 1;cactus_sprite[3][21][6] = 1;cactus_sprite[3][21][7] = 1;cactus_sprite[3][21][8] = 1;cactus_sprite[3][21][9] = 1;cactus_sprite[3][21][10] = 1;cactus_sprite[3][21][11] = 1;cactus_sprite[3][21][12] = 1;cactus_sprite[3][21][13] = 1;cactus_sprite[3][21][14] = 1;cactus_sprite[3][21][15] = 1;cactus_sprite[3][21][16] = 1;cactus_sprite[3][21][17] = 1;cactus_sprite[3][21][18] = 1;cactus_sprite[3][21][19] = 1;cactus_sprite[3][21][20] = 1;cactus_sprite[3][21][21] = 1;cactus_sprite[3][21][22] = 1;cactus_sprite[3][21][23] = 1;cactus_sprite[3][21][24] = 1;cactus_sprite[3][21][25] = 1;cactus_sprite[3][21][26] = 1;cactus_sprite[3][21][27] = 1;cactus_sprite[3][21][28] = 1;cactus_sprite[3][21][29] = 1;cactus_sprite[3][21][30] = 1;cactus_sprite[3][21][31] = 1;cactus_sprite[3][21][32] = 1;cactus_sprite[3][21][33] = 1;cactus_sprite[3][21][34] = 1;cactus_sprite[3][21][35] = 1;cactus_sprite[3][21][36] = 1;cactus_sprite[3][21][37] = 1;cactus_sprite[3][21][38] = 1;cactus_sprite[3][21][39] = 1;cactus_sprite[3][21][40] = 1;cactus_sprite[3][21][41] = 1;cactus_sprite[3][21][42] = 1;cactus_sprite[3][21][43] = 1;cactus_sprite[3][21][44] = 1;cactus_sprite[3][21][45] = 1;cactus_sprite[3][21][46] = 1;cactus_sprite[3][21][47] = 1;cactus_sprite[3][21][48] = 1;cactus_sprite[3][21][49] = 1;cactus_sprite[3][21][50] = 1;cactus_sprite[3][21][51] = 1;cactus_sprite[3][21][52] = 1;cactus_sprite[3][21][53] = 1;cactus_sprite[3][21][54] = 1;cactus_sprite[3][21][55] = 1;cactus_sprite[3][21][56] = 1;cactus_sprite[3][21][57] = 1;cactus_sprite[3][21][58] = 1;cactus_sprite[3][21][59] = 1;cactus_sprite[3][21][60] = 1;cactus_sprite[3][21][61] = 1;cactus_sprite[3][21][62] = 1;cactus_sprite[3][21][63] = 1;cactus_sprite[3][21][64] = 1;cactus_sprite[3][21][65] = 1;cactus_sprite[3][21][66] = 1;cactus_sprite[3][21][67] = 1;cactus_sprite[3][21][68] = 1;cactus_sprite[3][21][69] = 1;cactus_sprite[3][21][70] = 1;cactus_sprite[3][21][71] = 1;cactus_sprite[3][21][72] = 1;cactus_sprite[3][21][73] = 1;cactus_sprite[3][21][74] = 1;cactus_sprite[3][21][75] = 1;cactus_sprite[3][21][76] = 1;cactus_sprite[3][21][77] = 1;cactus_sprite[3][21][78] = 1;cactus_sprite[3][21][79] = 1;cactus_sprite[3][21][80] = 1;cactus_sprite[3][21][81] = 1;cactus_sprite[3][21][82] = 1;cactus_sprite[3][21][83] = 1;cactus_sprite[3][21][84] = 1;cactus_sprite[3][21][85] = 1;cactus_sprite[3][21][86] = 1;cactus_sprite[3][21][87] = 1;cactus_sprite[3][21][88] = 1;cactus_sprite[3][21][89] = 1;cactus_sprite[3][21][90] = 1;cactus_sprite[3][21][91] = 1;cactus_sprite[3][21][92] = 1;cactus_sprite[3][21][93] = 1;cactus_sprite[3][21][94] = 1;cactus_sprite[3][21][95] = 1;cactus_sprite[3][21][96] = 1;cactus_sprite[3][21][97] = 1;cactus_sprite[3][21][98] = 1;cactus_sprite[3][21][99] = 1;cactus_sprite[3][22][6] = 1;cactus_sprite[3][22][7] = 1;cactus_sprite[3][22][8] = 1;cactus_sprite[3][22][9] = 1;cactus_sprite[3][22][10] = 1;cactus_sprite[3][22][11] = 1;cactus_sprite[3][22][12] = 1;cactus_sprite[3][22][13] = 1;cactus_sprite[3][22][14] = 1;cactus_sprite[3][22][15] = 1;cactus_sprite[3][22][16] = 1;cactus_sprite[3][22][17] = 1;cactus_sprite[3][22][18] = 1;cactus_sprite[3][22][19] = 1;cactus_sprite[3][22][20] = 1;cactus_sprite[3][22][21] = 1;cactus_sprite[3][22][22] = 1;cactus_sprite[3][22][23] = 1;cactus_sprite[3][22][24] = 1;cactus_sprite[3][22][25] = 1;cactus_sprite[3][22][26] = 1;cactus_sprite[3][22][27] = 1;cactus_sprite[3][22][28] = 1;cactus_sprite[3][22][29] = 1;cactus_sprite[3][22][30] = 1;cactus_sprite[3][22][31] = 1;cactus_sprite[3][22][32] = 1;cactus_sprite[3][22][33] = 1;cactus_sprite[3][22][34] = 1;cactus_sprite[3][22][35] = 1;cactus_sprite[3][22][36] = 1;cactus_sprite[3][22][37] = 1;cactus_sprite[3][22][38] = 1;cactus_sprite[3][22][39] = 1;cactus_sprite[3][22][40] = 1;cactus_sprite[3][22][41] = 1;cactus_sprite[3][22][42] = 1;cactus_sprite[3][22][43] = 1;cactus_sprite[3][22][44] = 1;cactus_sprite[3][22][45] = 1;cactus_sprite[3][22][46] = 1;cactus_sprite[3][22][47] = 1;cactus_sprite[3][22][48] = 1;cactus_sprite[3][22][49] = 1;cactus_sprite[3][22][50] = 1;cactus_sprite[3][22][51] = 1;cactus_sprite[3][22][52] = 1;cactus_sprite[3][22][53] = 1;cactus_sprite[3][22][54] = 1;cactus_sprite[3][22][55] = 1;cactus_sprite[3][22][56] = 1;cactus_sprite[3][22][57] = 1;cactus_sprite[3][22][58] = 1;cactus_sprite[3][22][59] = 1;cactus_sprite[3][22][60] = 1;cactus_sprite[3][22][61] = 1;cactus_sprite[3][22][62] = 1;cactus_sprite[3][22][63] = 1;cactus_sprite[3][22][64] = 1;cactus_sprite[3][22][65] = 1;cactus_sprite[3][22][66] = 1;cactus_sprite[3][22][67] = 1;cactus_sprite[3][22][68] = 1;cactus_sprite[3][22][69] = 1;cactus_sprite[3][22][70] = 1;cactus_sprite[3][22][71] = 1;cactus_sprite[3][22][72] = 1;cactus_sprite[3][22][73] = 1;cactus_sprite[3][22][74] = 1;cactus_sprite[3][22][75] = 1;cactus_sprite[3][22][76] = 1;cactus_sprite[3][22][77] = 1;cactus_sprite[3][22][78] = 1;cactus_sprite[3][22][79] = 1;cactus_sprite[3][22][80] = 1;cactus_sprite[3][22][81] = 1;cactus_sprite[3][22][82] = 1;cactus_sprite[3][22][83] = 1;cactus_sprite[3][22][84] = 1;cactus_sprite[3][22][85] = 1;cactus_sprite[3][22][86] = 1;cactus_sprite[3][22][87] = 1;cactus_sprite[3][22][88] = 1;cactus_sprite[3][22][89] = 1;cactus_sprite[3][22][90] = 1;cactus_sprite[3][22][91] = 1;cactus_sprite[3][22][92] = 1;cactus_sprite[3][22][93] = 1;cactus_sprite[3][22][94] = 1;cactus_sprite[3][22][95] = 1;cactus_sprite[3][22][96] = 1;cactus_sprite[3][22][97] = 1;cactus_sprite[3][22][98] = 1;cactus_sprite[3][22][99] = 1;cactus_sprite[3][23][6] = 1;cactus_sprite[3][23][7] = 1;cactus_sprite[3][23][8] = 1;cactus_sprite[3][23][9] = 1;cactus_sprite[3][23][10] = 1;cactus_sprite[3][23][11] = 1;cactus_sprite[3][23][12] = 1;cactus_sprite[3][23][13] = 1;cactus_sprite[3][23][14] = 1;cactus_sprite[3][23][15] = 1;cactus_sprite[3][23][16] = 1;cactus_sprite[3][23][17] = 1;cactus_sprite[3][23][18] = 1;cactus_sprite[3][23][19] = 1;cactus_sprite[3][23][20] = 1;cactus_sprite[3][23][21] = 1;cactus_sprite[3][23][22] = 1;cactus_sprite[3][23][23] = 1;cactus_sprite[3][23][24] = 1;cactus_sprite[3][23][25] = 1;cactus_sprite[3][23][26] = 1;cactus_sprite[3][23][27] = 1;cactus_sprite[3][23][28] = 1;cactus_sprite[3][23][29] = 1;cactus_sprite[3][23][30] = 1;cactus_sprite[3][23][31] = 1;cactus_sprite[3][23][32] = 1;cactus_sprite[3][23][33] = 1;cactus_sprite[3][23][34] = 1;cactus_sprite[3][23][35] = 1;cactus_sprite[3][23][36] = 1;cactus_sprite[3][23][37] = 1;cactus_sprite[3][23][38] = 1;cactus_sprite[3][23][39] = 1;cactus_sprite[3][23][40] = 1;cactus_sprite[3][23][41] = 1;cactus_sprite[3][23][42] = 1;cactus_sprite[3][23][43] = 1;cactus_sprite[3][23][44] = 1;cactus_sprite[3][23][45] = 1;cactus_sprite[3][23][46] = 1;cactus_sprite[3][23][47] = 1;cactus_sprite[3][23][48] = 1;cactus_sprite[3][23][49] = 1;cactus_sprite[3][23][50] = 1;cactus_sprite[3][23][51] = 1;cactus_sprite[3][23][52] = 1;cactus_sprite[3][23][53] = 1;cactus_sprite[3][23][54] = 1;cactus_sprite[3][23][55] = 1;cactus_sprite[3][23][56] = 1;cactus_sprite[3][23][57] = 1;cactus_sprite[3][23][58] = 1;cactus_sprite[3][23][59] = 1;cactus_sprite[3][23][60] = 1;cactus_sprite[3][23][61] = 1;cactus_sprite[3][23][62] = 1;cactus_sprite[3][23][63] = 1;cactus_sprite[3][23][64] = 1;cactus_sprite[3][23][65] = 1;cactus_sprite[3][23][66] = 1;cactus_sprite[3][23][67] = 1;cactus_sprite[3][23][68] = 1;cactus_sprite[3][23][69] = 1;cactus_sprite[3][23][70] = 1;cactus_sprite[3][23][71] = 1;cactus_sprite[3][23][72] = 1;cactus_sprite[3][23][73] = 1;cactus_sprite[3][23][74] = 1;cactus_sprite[3][23][75] = 1;cactus_sprite[3][23][76] = 1;cactus_sprite[3][23][77] = 1;cactus_sprite[3][23][78] = 1;cactus_sprite[3][23][79] = 1;cactus_sprite[3][23][80] = 1;cactus_sprite[3][23][81] = 1;cactus_sprite[3][23][82] = 1;cactus_sprite[3][23][83] = 1;cactus_sprite[3][23][84] = 1;cactus_sprite[3][23][85] = 1;cactus_sprite[3][23][86] = 1;cactus_sprite[3][23][87] = 1;cactus_sprite[3][23][88] = 1;cactus_sprite[3][23][89] = 1;cactus_sprite[3][23][90] = 1;cactus_sprite[3][23][91] = 1;cactus_sprite[3][23][92] = 1;cactus_sprite[3][23][93] = 1;cactus_sprite[3][23][94] = 1;cactus_sprite[3][23][95] = 1;cactus_sprite[3][23][96] = 1;cactus_sprite[3][23][97] = 1;cactus_sprite[3][23][98] = 1;cactus_sprite[3][23][99] = 1;cactus_sprite[3][24][6] = 1;cactus_sprite[3][24][7] = 1;cactus_sprite[3][24][8] = 1;cactus_sprite[3][24][9] = 1;cactus_sprite[3][24][10] = 1;cactus_sprite[3][24][11] = 1;cactus_sprite[3][24][12] = 1;cactus_sprite[3][24][13] = 1;cactus_sprite[3][24][14] = 1;cactus_sprite[3][24][15] = 1;cactus_sprite[3][24][16] = 1;cactus_sprite[3][24][17] = 1;cactus_sprite[3][24][18] = 1;cactus_sprite[3][24][19] = 1;cactus_sprite[3][24][20] = 1;cactus_sprite[3][24][21] = 1;cactus_sprite[3][24][22] = 1;cactus_sprite[3][24][23] = 1;cactus_sprite[3][24][24] = 1;cactus_sprite[3][24][25] = 1;cactus_sprite[3][24][26] = 1;cactus_sprite[3][24][27] = 1;cactus_sprite[3][24][28] = 1;cactus_sprite[3][24][29] = 1;cactus_sprite[3][24][30] = 1;cactus_sprite[3][24][31] = 1;cactus_sprite[3][24][32] = 1;cactus_sprite[3][24][33] = 1;cactus_sprite[3][24][34] = 1;cactus_sprite[3][24][35] = 1;cactus_sprite[3][24][36] = 1;cactus_sprite[3][24][37] = 1;cactus_sprite[3][24][38] = 1;cactus_sprite[3][24][39] = 1;cactus_sprite[3][24][40] = 1;cactus_sprite[3][24][41] = 1;cactus_sprite[3][24][42] = 1;cactus_sprite[3][24][43] = 1;cactus_sprite[3][24][44] = 1;cactus_sprite[3][24][45] = 1;cactus_sprite[3][24][46] = 1;cactus_sprite[3][24][47] = 1;cactus_sprite[3][24][48] = 1;cactus_sprite[3][24][49] = 1;cactus_sprite[3][24][50] = 1;cactus_sprite[3][24][51] = 1;cactus_sprite[3][24][52] = 1;cactus_sprite[3][24][53] = 1;cactus_sprite[3][24][54] = 1;cactus_sprite[3][24][55] = 1;cactus_sprite[3][24][56] = 1;cactus_sprite[3][24][57] = 1;cactus_sprite[3][24][58] = 1;cactus_sprite[3][24][59] = 1;cactus_sprite[3][24][60] = 1;cactus_sprite[3][24][61] = 1;cactus_sprite[3][24][62] = 1;cactus_sprite[3][24][63] = 1;cactus_sprite[3][24][64] = 1;cactus_sprite[3][24][65] = 1;cactus_sprite[3][24][66] = 1;cactus_sprite[3][24][67] = 1;cactus_sprite[3][24][68] = 1;cactus_sprite[3][24][69] = 1;cactus_sprite[3][24][70] = 1;cactus_sprite[3][24][71] = 1;cactus_sprite[3][24][72] = 1;cactus_sprite[3][24][73] = 1;cactus_sprite[3][24][74] = 1;cactus_sprite[3][24][75] = 1;cactus_sprite[3][24][76] = 1;cactus_sprite[3][24][77] = 1;cactus_sprite[3][24][78] = 1;cactus_sprite[3][24][79] = 1;cactus_sprite[3][24][80] = 1;cactus_sprite[3][24][81] = 1;cactus_sprite[3][24][82] = 1;cactus_sprite[3][24][83] = 1;cactus_sprite[3][24][84] = 1;cactus_sprite[3][24][85] = 1;cactus_sprite[3][24][86] = 1;cactus_sprite[3][24][87] = 1;cactus_sprite[3][24][88] = 1;cactus_sprite[3][24][89] = 1;cactus_sprite[3][24][90] = 1;cactus_sprite[3][24][91] = 1;cactus_sprite[3][24][92] = 1;cactus_sprite[3][24][93] = 1;cactus_sprite[3][24][94] = 1;cactus_sprite[3][24][95] = 1;cactus_sprite[3][24][96] = 1;cactus_sprite[3][24][97] = 1;cactus_sprite[3][24][98] = 1;cactus_sprite[3][24][99] = 1;cactus_sprite[3][25][6] = 1;cactus_sprite[3][25][7] = 1;cactus_sprite[3][25][8] = 1;cactus_sprite[3][25][9] = 1;cactus_sprite[3][25][10] = 1;cactus_sprite[3][25][11] = 1;cactus_sprite[3][25][12] = 1;cactus_sprite[3][25][13] = 1;cactus_sprite[3][25][14] = 1;cactus_sprite[3][25][15] = 1;cactus_sprite[3][25][16] = 1;cactus_sprite[3][25][17] = 1;cactus_sprite[3][25][18] = 1;cactus_sprite[3][25][19] = 1;cactus_sprite[3][25][20] = 1;cactus_sprite[3][25][21] = 1;cactus_sprite[3][25][22] = 1;cactus_sprite[3][25][23] = 1;cactus_sprite[3][25][24] = 1;cactus_sprite[3][25][25] = 1;cactus_sprite[3][25][26] = 1;cactus_sprite[3][25][27] = 1;cactus_sprite[3][25][28] = 1;cactus_sprite[3][25][29] = 1;cactus_sprite[3][25][30] = 1;cactus_sprite[3][25][31] = 1;cactus_sprite[3][25][32] = 1;cactus_sprite[3][25][33] = 1;cactus_sprite[3][25][34] = 1;cactus_sprite[3][25][35] = 1;cactus_sprite[3][25][36] = 1;cactus_sprite[3][25][37] = 1;cactus_sprite[3][25][38] = 1;cactus_sprite[3][25][39] = 1;cactus_sprite[3][25][40] = 1;cactus_sprite[3][25][41] = 1;cactus_sprite[3][25][42] = 1;cactus_sprite[3][25][43] = 1;cactus_sprite[3][25][44] = 1;cactus_sprite[3][25][45] = 1;cactus_sprite[3][25][46] = 1;cactus_sprite[3][25][47] = 1;cactus_sprite[3][25][48] = 1;cactus_sprite[3][25][49] = 1;cactus_sprite[3][25][50] = 1;cactus_sprite[3][25][51] = 1;cactus_sprite[3][25][52] = 1;cactus_sprite[3][25][53] = 1;cactus_sprite[3][25][54] = 1;cactus_sprite[3][25][55] = 1;cactus_sprite[3][25][56] = 1;cactus_sprite[3][25][57] = 1;cactus_sprite[3][25][58] = 1;cactus_sprite[3][25][59] = 1;cactus_sprite[3][25][60] = 1;cactus_sprite[3][25][61] = 1;cactus_sprite[3][25][62] = 1;cactus_sprite[3][25][63] = 1;cactus_sprite[3][25][64] = 1;cactus_sprite[3][25][65] = 1;cactus_sprite[3][25][66] = 1;cactus_sprite[3][25][67] = 1;cactus_sprite[3][25][68] = 1;cactus_sprite[3][25][69] = 1;cactus_sprite[3][25][70] = 1;cactus_sprite[3][25][71] = 1;cactus_sprite[3][25][72] = 1;cactus_sprite[3][25][73] = 1;cactus_sprite[3][25][74] = 1;cactus_sprite[3][25][75] = 1;cactus_sprite[3][25][76] = 1;cactus_sprite[3][25][77] = 1;cactus_sprite[3][25][78] = 1;cactus_sprite[3][25][79] = 1;cactus_sprite[3][25][80] = 1;cactus_sprite[3][25][81] = 1;cactus_sprite[3][25][82] = 1;cactus_sprite[3][25][83] = 1;cactus_sprite[3][25][84] = 1;cactus_sprite[3][25][85] = 1;cactus_sprite[3][25][86] = 1;cactus_sprite[3][25][87] = 1;cactus_sprite[3][25][88] = 1;cactus_sprite[3][25][89] = 1;cactus_sprite[3][25][90] = 1;cactus_sprite[3][25][91] = 1;cactus_sprite[3][25][92] = 1;cactus_sprite[3][25][93] = 1;cactus_sprite[3][25][94] = 1;cactus_sprite[3][25][95] = 1;cactus_sprite[3][25][96] = 1;cactus_sprite[3][25][97] = 1;cactus_sprite[3][25][98] = 1;cactus_sprite[3][25][99] = 1;cactus_sprite[3][26][6] = 1;cactus_sprite[3][26][7] = 1;cactus_sprite[3][26][8] = 1;cactus_sprite[3][26][9] = 1;cactus_sprite[3][26][10] = 1;cactus_sprite[3][26][11] = 1;cactus_sprite[3][26][12] = 1;cactus_sprite[3][26][13] = 1;cactus_sprite[3][26][14] = 1;cactus_sprite[3][26][15] = 1;cactus_sprite[3][26][16] = 1;cactus_sprite[3][26][17] = 1;cactus_sprite[3][26][18] = 1;cactus_sprite[3][26][19] = 1;cactus_sprite[3][26][20] = 1;cactus_sprite[3][26][21] = 1;cactus_sprite[3][26][22] = 1;cactus_sprite[3][26][23] = 1;cactus_sprite[3][26][24] = 1;cactus_sprite[3][26][25] = 1;cactus_sprite[3][26][26] = 1;cactus_sprite[3][26][27] = 1;cactus_sprite[3][26][28] = 1;cactus_sprite[3][26][29] = 1;cactus_sprite[3][26][30] = 1;cactus_sprite[3][26][31] = 1;cactus_sprite[3][26][32] = 1;cactus_sprite[3][26][33] = 1;cactus_sprite[3][26][34] = 1;cactus_sprite[3][26][35] = 1;cactus_sprite[3][26][36] = 1;cactus_sprite[3][26][37] = 1;cactus_sprite[3][26][38] = 1;cactus_sprite[3][26][39] = 1;cactus_sprite[3][26][40] = 1;cactus_sprite[3][26][41] = 1;cactus_sprite[3][26][42] = 1;cactus_sprite[3][26][43] = 1;cactus_sprite[3][26][44] = 1;cactus_sprite[3][26][45] = 1;cactus_sprite[3][26][46] = 1;cactus_sprite[3][26][47] = 1;cactus_sprite[3][26][48] = 1;cactus_sprite[3][26][49] = 1;cactus_sprite[3][26][50] = 1;cactus_sprite[3][26][51] = 1;cactus_sprite[3][26][52] = 1;cactus_sprite[3][26][53] = 1;cactus_sprite[3][26][54] = 1;cactus_sprite[3][26][55] = 1;cactus_sprite[3][26][56] = 1;cactus_sprite[3][26][57] = 1;cactus_sprite[3][26][58] = 1;cactus_sprite[3][26][59] = 1;cactus_sprite[3][26][60] = 1;cactus_sprite[3][26][61] = 1;cactus_sprite[3][26][62] = 1;cactus_sprite[3][26][63] = 1;cactus_sprite[3][26][64] = 1;cactus_sprite[3][26][65] = 1;cactus_sprite[3][26][66] = 1;cactus_sprite[3][26][67] = 1;cactus_sprite[3][26][68] = 1;cactus_sprite[3][26][69] = 1;cactus_sprite[3][26][70] = 1;cactus_sprite[3][26][71] = 1;cactus_sprite[3][26][72] = 1;cactus_sprite[3][26][73] = 1;cactus_sprite[3][26][74] = 1;cactus_sprite[3][26][75] = 1;cactus_sprite[3][26][76] = 1;cactus_sprite[3][26][77] = 1;cactus_sprite[3][26][78] = 1;cactus_sprite[3][26][79] = 1;cactus_sprite[3][26][80] = 1;cactus_sprite[3][26][81] = 1;cactus_sprite[3][26][82] = 1;cactus_sprite[3][26][83] = 1;cactus_sprite[3][26][84] = 1;cactus_sprite[3][26][85] = 1;cactus_sprite[3][26][86] = 1;cactus_sprite[3][26][87] = 1;cactus_sprite[3][26][88] = 1;cactus_sprite[3][26][89] = 1;cactus_sprite[3][26][90] = 1;cactus_sprite[3][26][91] = 1;cactus_sprite[3][26][92] = 1;cactus_sprite[3][26][93] = 1;cactus_sprite[3][26][94] = 1;cactus_sprite[3][26][95] = 1;cactus_sprite[3][26][96] = 1;cactus_sprite[3][26][97] = 1;cactus_sprite[3][26][98] = 1;cactus_sprite[3][26][99] = 1;cactus_sprite[3][27][6] = 1;cactus_sprite[3][27][7] = 1;cactus_sprite[3][27][8] = 1;cactus_sprite[3][27][9] = 1;cactus_sprite[3][27][10] = 1;cactus_sprite[3][27][11] = 1;cactus_sprite[3][27][12] = 1;cactus_sprite[3][27][13] = 1;cactus_sprite[3][27][14] = 1;cactus_sprite[3][27][15] = 1;cactus_sprite[3][27][16] = 1;cactus_sprite[3][27][17] = 1;cactus_sprite[3][27][18] = 1;cactus_sprite[3][27][19] = 1;cactus_sprite[3][27][20] = 1;cactus_sprite[3][27][21] = 1;cactus_sprite[3][27][22] = 1;cactus_sprite[3][27][23] = 1;cactus_sprite[3][27][24] = 1;cactus_sprite[3][27][25] = 1;cactus_sprite[3][27][26] = 1;cactus_sprite[3][27][27] = 1;cactus_sprite[3][27][28] = 1;cactus_sprite[3][27][29] = 1;cactus_sprite[3][27][30] = 1;cactus_sprite[3][27][31] = 1;cactus_sprite[3][27][32] = 1;cactus_sprite[3][27][33] = 1;cactus_sprite[3][27][34] = 1;cactus_sprite[3][27][35] = 1;cactus_sprite[3][27][36] = 1;cactus_sprite[3][27][37] = 1;cactus_sprite[3][27][38] = 1;cactus_sprite[3][27][39] = 1;cactus_sprite[3][27][40] = 1;cactus_sprite[3][27][41] = 1;cactus_sprite[3][27][42] = 1;cactus_sprite[3][27][43] = 1;cactus_sprite[3][27][44] = 1;cactus_sprite[3][27][45] = 1;cactus_sprite[3][27][46] = 1;cactus_sprite[3][27][47] = 1;cactus_sprite[3][27][48] = 1;cactus_sprite[3][27][49] = 1;cactus_sprite[3][27][50] = 1;cactus_sprite[3][27][51] = 1;cactus_sprite[3][27][52] = 1;cactus_sprite[3][27][53] = 1;cactus_sprite[3][27][54] = 1;cactus_sprite[3][27][55] = 1;cactus_sprite[3][27][56] = 1;cactus_sprite[3][27][57] = 1;cactus_sprite[3][27][58] = 1;cactus_sprite[3][27][59] = 1;cactus_sprite[3][27][60] = 1;cactus_sprite[3][27][61] = 1;cactus_sprite[3][27][62] = 1;cactus_sprite[3][27][63] = 1;cactus_sprite[3][27][64] = 1;cactus_sprite[3][27][65] = 1;cactus_sprite[3][27][66] = 1;cactus_sprite[3][27][67] = 1;cactus_sprite[3][27][68] = 1;cactus_sprite[3][27][69] = 1;cactus_sprite[3][27][70] = 1;cactus_sprite[3][27][71] = 1;cactus_sprite[3][27][72] = 1;cactus_sprite[3][27][73] = 1;cactus_sprite[3][27][74] = 1;cactus_sprite[3][27][75] = 1;cactus_sprite[3][27][76] = 1;cactus_sprite[3][27][77] = 1;cactus_sprite[3][27][78] = 1;cactus_sprite[3][27][79] = 1;cactus_sprite[3][27][80] = 1;cactus_sprite[3][27][81] = 1;cactus_sprite[3][27][82] = 1;cactus_sprite[3][27][83] = 1;cactus_sprite[3][27][84] = 1;cactus_sprite[3][27][85] = 1;cactus_sprite[3][27][86] = 1;cactus_sprite[3][27][87] = 1;cactus_sprite[3][27][88] = 1;cactus_sprite[3][27][89] = 1;cactus_sprite[3][27][90] = 1;cactus_sprite[3][27][91] = 1;cactus_sprite[3][27][92] = 1;cactus_sprite[3][27][93] = 1;cactus_sprite[3][27][94] = 1;cactus_sprite[3][27][95] = 1;cactus_sprite[3][27][96] = 1;cactus_sprite[3][27][97] = 1;cactus_sprite[3][27][98] = 1;cactus_sprite[3][27][99] = 1;cactus_sprite[3][28][6] = 1;cactus_sprite[3][28][7] = 1;cactus_sprite[3][28][8] = 1;cactus_sprite[3][28][9] = 1;cactus_sprite[3][28][10] = 1;cactus_sprite[3][28][11] = 1;cactus_sprite[3][28][12] = 1;cactus_sprite[3][28][13] = 1;cactus_sprite[3][28][14] = 1;cactus_sprite[3][28][15] = 1;cactus_sprite[3][28][16] = 1;cactus_sprite[3][28][17] = 1;cactus_sprite[3][28][18] = 1;cactus_sprite[3][28][19] = 1;cactus_sprite[3][28][20] = 1;cactus_sprite[3][28][21] = 1;cactus_sprite[3][28][22] = 1;cactus_sprite[3][28][23] = 1;cactus_sprite[3][28][24] = 1;cactus_sprite[3][28][25] = 1;cactus_sprite[3][28][26] = 1;cactus_sprite[3][28][27] = 1;cactus_sprite[3][28][28] = 1;cactus_sprite[3][28][29] = 1;cactus_sprite[3][28][30] = 1;cactus_sprite[3][28][31] = 1;cactus_sprite[3][28][32] = 1;cactus_sprite[3][28][33] = 1;cactus_sprite[3][28][34] = 1;cactus_sprite[3][28][35] = 1;cactus_sprite[3][28][36] = 1;cactus_sprite[3][28][37] = 1;cactus_sprite[3][28][38] = 1;cactus_sprite[3][28][39] = 1;cactus_sprite[3][28][40] = 1;cactus_sprite[3][28][41] = 1;cactus_sprite[3][28][42] = 1;cactus_sprite[3][28][43] = 1;cactus_sprite[3][28][44] = 1;cactus_sprite[3][28][45] = 1;cactus_sprite[3][28][46] = 1;cactus_sprite[3][28][47] = 1;cactus_sprite[3][28][48] = 1;cactus_sprite[3][28][49] = 1;cactus_sprite[3][28][50] = 1;cactus_sprite[3][28][51] = 1;cactus_sprite[3][28][52] = 1;cactus_sprite[3][28][53] = 1;cactus_sprite[3][28][54] = 1;cactus_sprite[3][28][55] = 1;cactus_sprite[3][28][56] = 1;cactus_sprite[3][28][57] = 1;cactus_sprite[3][28][58] = 1;cactus_sprite[3][28][59] = 1;cactus_sprite[3][28][60] = 1;cactus_sprite[3][28][61] = 1;cactus_sprite[3][28][62] = 1;cactus_sprite[3][28][63] = 1;cactus_sprite[3][28][64] = 1;cactus_sprite[3][28][65] = 1;cactus_sprite[3][28][66] = 1;cactus_sprite[3][28][67] = 1;cactus_sprite[3][28][68] = 1;cactus_sprite[3][28][69] = 1;cactus_sprite[3][28][70] = 1;cactus_sprite[3][28][71] = 1;cactus_sprite[3][28][72] = 1;cactus_sprite[3][28][73] = 1;cactus_sprite[3][28][74] = 1;cactus_sprite[3][28][75] = 1;cactus_sprite[3][28][76] = 1;cactus_sprite[3][28][77] = 1;cactus_sprite[3][28][78] = 1;cactus_sprite[3][28][79] = 1;cactus_sprite[3][28][80] = 1;cactus_sprite[3][28][81] = 1;cactus_sprite[3][28][82] = 1;cactus_sprite[3][28][83] = 1;cactus_sprite[3][28][84] = 1;cactus_sprite[3][28][85] = 1;cactus_sprite[3][28][86] = 1;cactus_sprite[3][28][87] = 1;cactus_sprite[3][28][88] = 1;cactus_sprite[3][28][89] = 1;cactus_sprite[3][28][90] = 1;cactus_sprite[3][28][91] = 1;cactus_sprite[3][28][92] = 1;cactus_sprite[3][28][93] = 1;cactus_sprite[3][28][94] = 1;cactus_sprite[3][28][95] = 1;cactus_sprite[3][28][96] = 1;cactus_sprite[3][28][97] = 1;cactus_sprite[3][28][98] = 1;cactus_sprite[3][28][99] = 1;cactus_sprite[3][29][6] = 1;cactus_sprite[3][29][7] = 1;cactus_sprite[3][29][8] = 1;cactus_sprite[3][29][9] = 1;cactus_sprite[3][29][10] = 1;cactus_sprite[3][29][11] = 1;cactus_sprite[3][29][12] = 1;cactus_sprite[3][29][13] = 1;cactus_sprite[3][29][14] = 1;cactus_sprite[3][29][15] = 1;cactus_sprite[3][29][16] = 1;cactus_sprite[3][29][17] = 1;cactus_sprite[3][29][18] = 1;cactus_sprite[3][29][19] = 1;cactus_sprite[3][29][20] = 1;cactus_sprite[3][29][21] = 1;cactus_sprite[3][29][22] = 1;cactus_sprite[3][29][23] = 1;cactus_sprite[3][29][24] = 1;cactus_sprite[3][29][25] = 1;cactus_sprite[3][29][26] = 1;cactus_sprite[3][29][27] = 1;cactus_sprite[3][29][28] = 1;cactus_sprite[3][29][29] = 1;cactus_sprite[3][29][30] = 1;cactus_sprite[3][29][31] = 1;cactus_sprite[3][29][32] = 1;cactus_sprite[3][29][33] = 1;cactus_sprite[3][29][34] = 1;cactus_sprite[3][29][35] = 1;cactus_sprite[3][29][36] = 1;cactus_sprite[3][29][37] = 1;cactus_sprite[3][29][38] = 1;cactus_sprite[3][29][39] = 1;cactus_sprite[3][29][40] = 1;cactus_sprite[3][29][41] = 1;cactus_sprite[3][29][42] = 1;cactus_sprite[3][29][43] = 1;cactus_sprite[3][29][44] = 1;cactus_sprite[3][29][45] = 1;cactus_sprite[3][29][46] = 1;cactus_sprite[3][29][47] = 1;cactus_sprite[3][29][48] = 1;cactus_sprite[3][29][49] = 1;cactus_sprite[3][29][50] = 1;cactus_sprite[3][29][51] = 1;cactus_sprite[3][29][52] = 1;cactus_sprite[3][29][53] = 1;cactus_sprite[3][29][54] = 1;cactus_sprite[3][29][55] = 1;cactus_sprite[3][29][56] = 1;cactus_sprite[3][29][57] = 1;cactus_sprite[3][29][58] = 1;cactus_sprite[3][29][59] = 1;cactus_sprite[3][29][60] = 1;cactus_sprite[3][29][61] = 1;cactus_sprite[3][29][62] = 1;cactus_sprite[3][29][63] = 1;cactus_sprite[3][29][64] = 1;cactus_sprite[3][29][65] = 1;cactus_sprite[3][29][66] = 1;cactus_sprite[3][29][67] = 1;cactus_sprite[3][29][68] = 1;cactus_sprite[3][29][69] = 1;cactus_sprite[3][29][70] = 1;cactus_sprite[3][29][71] = 1;cactus_sprite[3][29][72] = 1;cactus_sprite[3][29][73] = 1;cactus_sprite[3][29][74] = 1;cactus_sprite[3][29][75] = 1;cactus_sprite[3][29][76] = 1;cactus_sprite[3][29][77] = 1;cactus_sprite[3][29][78] = 1;cactus_sprite[3][29][79] = 1;cactus_sprite[3][29][80] = 1;cactus_sprite[3][29][81] = 1;cactus_sprite[3][29][82] = 1;cactus_sprite[3][29][83] = 1;cactus_sprite[3][29][84] = 1;cactus_sprite[3][29][85] = 1;cactus_sprite[3][29][86] = 1;cactus_sprite[3][29][87] = 1;cactus_sprite[3][29][88] = 1;cactus_sprite[3][29][89] = 1;cactus_sprite[3][29][90] = 1;cactus_sprite[3][29][91] = 1;cactus_sprite[3][29][92] = 1;cactus_sprite[3][29][93] = 1;cactus_sprite[3][29][94] = 1;cactus_sprite[3][29][95] = 1;cactus_sprite[3][29][96] = 1;cactus_sprite[3][29][97] = 1;cactus_sprite[3][29][98] = 1;cactus_sprite[3][29][99] = 1;cactus_sprite[3][30][8] = 1;cactus_sprite[3][30][9] = 1;cactus_sprite[3][30][10] = 1;cactus_sprite[3][30][11] = 1;cactus_sprite[3][30][12] = 1;cactus_sprite[3][30][13] = 1;cactus_sprite[3][30][14] = 1;cactus_sprite[3][30][15] = 1;cactus_sprite[3][30][16] = 1;cactus_sprite[3][30][17] = 1;cactus_sprite[3][30][18] = 1;cactus_sprite[3][30][19] = 1;cactus_sprite[3][30][20] = 1;cactus_sprite[3][30][21] = 1;cactus_sprite[3][30][22] = 1;cactus_sprite[3][30][23] = 1;cactus_sprite[3][30][24] = 1;cactus_sprite[3][30][25] = 1;cactus_sprite[3][30][26] = 1;cactus_sprite[3][30][27] = 1;cactus_sprite[3][30][28] = 1;cactus_sprite[3][30][29] = 1;cactus_sprite[3][30][30] = 1;cactus_sprite[3][30][31] = 1;cactus_sprite[3][30][32] = 1;cactus_sprite[3][30][33] = 1;cactus_sprite[3][30][34] = 1;cactus_sprite[3][30][35] = 1;cactus_sprite[3][30][36] = 1;cactus_sprite[3][30][37] = 1;cactus_sprite[3][30][38] = 1;cactus_sprite[3][30][39] = 1;cactus_sprite[3][30][40] = 1;cactus_sprite[3][30][41] = 1;cactus_sprite[3][30][42] = 1;cactus_sprite[3][30][43] = 1;cactus_sprite[3][30][44] = 1;cactus_sprite[3][30][45] = 1;cactus_sprite[3][30][46] = 1;cactus_sprite[3][30][47] = 1;cactus_sprite[3][30][48] = 1;cactus_sprite[3][30][49] = 1;cactus_sprite[3][30][50] = 1;cactus_sprite[3][30][51] = 1;cactus_sprite[3][30][52] = 1;cactus_sprite[3][30][53] = 1;cactus_sprite[3][30][54] = 1;cactus_sprite[3][30][55] = 1;cactus_sprite[3][30][56] = 1;cactus_sprite[3][30][57] = 1;cactus_sprite[3][30][58] = 1;cactus_sprite[3][30][59] = 1;cactus_sprite[3][30][60] = 1;cactus_sprite[3][30][61] = 1;cactus_sprite[3][30][62] = 1;cactus_sprite[3][30][63] = 1;cactus_sprite[3][30][64] = 1;cactus_sprite[3][30][65] = 1;cactus_sprite[3][30][66] = 1;cactus_sprite[3][30][67] = 1;cactus_sprite[3][30][68] = 1;cactus_sprite[3][30][69] = 1;cactus_sprite[3][30][70] = 1;cactus_sprite[3][30][71] = 1;cactus_sprite[3][30][72] = 1;cactus_sprite[3][30][73] = 1;cactus_sprite[3][30][74] = 1;cactus_sprite[3][30][75] = 1;cactus_sprite[3][30][76] = 1;cactus_sprite[3][30][77] = 1;cactus_sprite[3][30][78] = 1;cactus_sprite[3][30][79] = 1;cactus_sprite[3][30][80] = 1;cactus_sprite[3][30][81] = 1;cactus_sprite[3][30][82] = 1;cactus_sprite[3][30][83] = 1;cactus_sprite[3][30][84] = 1;cactus_sprite[3][30][85] = 1;cactus_sprite[3][30][86] = 1;cactus_sprite[3][30][87] = 1;cactus_sprite[3][30][88] = 1;cactus_sprite[3][30][89] = 1;cactus_sprite[3][30][90] = 1;cactus_sprite[3][30][91] = 1;cactus_sprite[3][30][92] = 1;cactus_sprite[3][30][93] = 1;cactus_sprite[3][30][94] = 1;cactus_sprite[3][30][95] = 1;cactus_sprite[3][30][96] = 1;cactus_sprite[3][30][97] = 1;cactus_sprite[3][30][98] = 1;cactus_sprite[3][30][99] = 1;cactus_sprite[3][31][8] = 1;cactus_sprite[3][31][9] = 1;cactus_sprite[3][31][10] = 1;cactus_sprite[3][31][11] = 1;cactus_sprite[3][31][12] = 1;cactus_sprite[3][31][13] = 1;cactus_sprite[3][31][14] = 1;cactus_sprite[3][31][15] = 1;cactus_sprite[3][31][16] = 1;cactus_sprite[3][31][17] = 1;cactus_sprite[3][31][18] = 1;cactus_sprite[3][31][19] = 1;cactus_sprite[3][31][20] = 1;cactus_sprite[3][31][21] = 1;cactus_sprite[3][31][22] = 1;cactus_sprite[3][31][23] = 1;cactus_sprite[3][31][24] = 1;cactus_sprite[3][31][25] = 1;cactus_sprite[3][31][26] = 1;cactus_sprite[3][31][27] = 1;cactus_sprite[3][31][28] = 1;cactus_sprite[3][31][29] = 1;cactus_sprite[3][31][30] = 1;cactus_sprite[3][31][31] = 1;cactus_sprite[3][31][32] = 1;cactus_sprite[3][31][33] = 1;cactus_sprite[3][31][34] = 1;cactus_sprite[3][31][35] = 1;cactus_sprite[3][31][36] = 1;cactus_sprite[3][31][37] = 1;cactus_sprite[3][31][38] = 1;cactus_sprite[3][31][39] = 1;cactus_sprite[3][31][40] = 1;cactus_sprite[3][31][41] = 1;cactus_sprite[3][31][42] = 1;cactus_sprite[3][31][43] = 1;cactus_sprite[3][31][44] = 1;cactus_sprite[3][31][45] = 1;cactus_sprite[3][31][46] = 1;cactus_sprite[3][31][47] = 1;cactus_sprite[3][31][48] = 1;cactus_sprite[3][31][49] = 1;cactus_sprite[3][31][50] = 1;cactus_sprite[3][31][51] = 1;cactus_sprite[3][31][52] = 1;cactus_sprite[3][31][53] = 1;cactus_sprite[3][31][54] = 1;cactus_sprite[3][31][55] = 1;cactus_sprite[3][31][56] = 1;cactus_sprite[3][31][57] = 1;cactus_sprite[3][31][58] = 1;cactus_sprite[3][31][59] = 1;cactus_sprite[3][31][60] = 1;cactus_sprite[3][31][61] = 1;cactus_sprite[3][31][62] = 1;cactus_sprite[3][31][63] = 1;cactus_sprite[3][31][64] = 1;cactus_sprite[3][31][65] = 1;cactus_sprite[3][31][66] = 1;cactus_sprite[3][31][67] = 1;cactus_sprite[3][31][68] = 1;cactus_sprite[3][31][69] = 1;cactus_sprite[3][31][70] = 1;cactus_sprite[3][31][71] = 1;cactus_sprite[3][31][72] = 1;cactus_sprite[3][31][73] = 1;cactus_sprite[3][31][74] = 1;cactus_sprite[3][31][75] = 1;cactus_sprite[3][31][76] = 1;cactus_sprite[3][31][77] = 1;cactus_sprite[3][31][78] = 1;cactus_sprite[3][31][79] = 1;cactus_sprite[3][31][80] = 1;cactus_sprite[3][31][81] = 1;cactus_sprite[3][31][82] = 1;cactus_sprite[3][31][83] = 1;cactus_sprite[3][31][84] = 1;cactus_sprite[3][31][85] = 1;cactus_sprite[3][31][86] = 1;cactus_sprite[3][31][87] = 1;cactus_sprite[3][31][88] = 1;cactus_sprite[3][31][89] = 1;cactus_sprite[3][31][90] = 1;cactus_sprite[3][31][91] = 1;cactus_sprite[3][31][92] = 1;cactus_sprite[3][31][93] = 1;cactus_sprite[3][31][94] = 1;cactus_sprite[3][31][95] = 1;cactus_sprite[3][31][96] = 1;cactus_sprite[3][31][97] = 1;cactus_sprite[3][31][98] = 1;cactus_sprite[3][31][99] = 1;cactus_sprite[3][32][60] = 1;cactus_sprite[3][32][61] = 1;cactus_sprite[3][32][62] = 1;cactus_sprite[3][32][63] = 1;cactus_sprite[3][32][64] = 1;cactus_sprite[3][32][65] = 1;cactus_sprite[3][33][60] = 1;cactus_sprite[3][33][61] = 1;cactus_sprite[3][33][62] = 1;cactus_sprite[3][33][63] = 1;cactus_sprite[3][33][64] = 1;cactus_sprite[3][33][65] = 1;cactus_sprite[3][34][60] = 1;cactus_sprite[3][34][61] = 1;cactus_sprite[3][34][62] = 1;cactus_sprite[3][34][63] = 1;cactus_sprite[3][34][64] = 1;cactus_sprite[3][34][65] = 1;cactus_sprite[3][35][60] = 1;cactus_sprite[3][35][61] = 1;cactus_sprite[3][35][62] = 1;cactus_sprite[3][35][63] = 1;cactus_sprite[3][35][64] = 1;cactus_sprite[3][35][65] = 1;cactus_sprite[3][36][60] = 1;cactus_sprite[3][36][61] = 1;cactus_sprite[3][36][62] = 1;cactus_sprite[3][36][63] = 1;cactus_sprite[3][36][64] = 1;cactus_sprite[3][36][65] = 1;cactus_sprite[3][37][60] = 1;cactus_sprite[3][37][61] = 1;cactus_sprite[3][37][62] = 1;cactus_sprite[3][37][63] = 1;cactus_sprite[3][37][64] = 1;cactus_sprite[3][37][65] = 1;cactus_sprite[3][38][30] = 1;cactus_sprite[3][38][31] = 1;cactus_sprite[3][38][32] = 1;cactus_sprite[3][38][33] = 1;cactus_sprite[3][38][34] = 1;cactus_sprite[3][38][35] = 1;cactus_sprite[3][38][36] = 1;cactus_sprite[3][38][37] = 1;cactus_sprite[3][38][38] = 1;cactus_sprite[3][38][39] = 1;cactus_sprite[3][38][40] = 1;cactus_sprite[3][38][41] = 1;cactus_sprite[3][38][42] = 1;cactus_sprite[3][38][43] = 1;cactus_sprite[3][38][44] = 1;cactus_sprite[3][38][45] = 1;cactus_sprite[3][38][46] = 1;cactus_sprite[3][38][47] = 1;cactus_sprite[3][38][48] = 1;cactus_sprite[3][38][49] = 1;cactus_sprite[3][38][50] = 1;cactus_sprite[3][38][51] = 1;cactus_sprite[3][38][52] = 1;cactus_sprite[3][38][53] = 1;cactus_sprite[3][38][54] = 1;cactus_sprite[3][38][55] = 1;cactus_sprite[3][38][56] = 1;cactus_sprite[3][38][57] = 1;cactus_sprite[3][38][58] = 1;cactus_sprite[3][38][59] = 1;cactus_sprite[3][38][60] = 1;cactus_sprite[3][38][61] = 1;cactus_sprite[3][38][62] = 1;cactus_sprite[3][38][63] = 1;cactus_sprite[3][38][64] = 1;cactus_sprite[3][38][65] = 1;cactus_sprite[3][39][30] = 1;cactus_sprite[3][39][31] = 1;cactus_sprite[3][39][32] = 1;cactus_sprite[3][39][33] = 1;cactus_sprite[3][39][34] = 1;cactus_sprite[3][39][35] = 1;cactus_sprite[3][39][36] = 1;cactus_sprite[3][39][37] = 1;cactus_sprite[3][39][38] = 1;cactus_sprite[3][39][39] = 1;cactus_sprite[3][39][40] = 1;cactus_sprite[3][39][41] = 1;cactus_sprite[3][39][42] = 1;cactus_sprite[3][39][43] = 1;cactus_sprite[3][39][44] = 1;cactus_sprite[3][39][45] = 1;cactus_sprite[3][39][46] = 1;cactus_sprite[3][39][47] = 1;cactus_sprite[3][39][48] = 1;cactus_sprite[3][39][49] = 1;cactus_sprite[3][39][50] = 1;cactus_sprite[3][39][51] = 1;cactus_sprite[3][39][52] = 1;cactus_sprite[3][39][53] = 1;cactus_sprite[3][39][54] = 1;cactus_sprite[3][39][55] = 1;cactus_sprite[3][39][56] = 1;cactus_sprite[3][39][57] = 1;cactus_sprite[3][39][58] = 1;cactus_sprite[3][39][59] = 1;cactus_sprite[3][39][60] = 1;cactus_sprite[3][39][61] = 1;cactus_sprite[3][39][62] = 1;cactus_sprite[3][39][63] = 1;cactus_sprite[3][39][64] = 1;cactus_sprite[3][39][65] = 1;cactus_sprite[3][40][28] = 1;cactus_sprite[3][40][29] = 1;cactus_sprite[3][40][30] = 1;cactus_sprite[3][40][31] = 1;cactus_sprite[3][40][32] = 1;cactus_sprite[3][40][33] = 1;cactus_sprite[3][40][34] = 1;cactus_sprite[3][40][35] = 1;cactus_sprite[3][40][36] = 1;cactus_sprite[3][40][37] = 1;cactus_sprite[3][40][38] = 1;cactus_sprite[3][40][39] = 1;cactus_sprite[3][40][40] = 1;cactus_sprite[3][40][41] = 1;cactus_sprite[3][40][42] = 1;cactus_sprite[3][40][43] = 1;cactus_sprite[3][40][44] = 1;cactus_sprite[3][40][45] = 1;cactus_sprite[3][40][46] = 1;cactus_sprite[3][40][47] = 1;cactus_sprite[3][40][48] = 1;cactus_sprite[3][40][49] = 1;cactus_sprite[3][40][50] = 1;cactus_sprite[3][40][51] = 1;cactus_sprite[3][40][52] = 1;cactus_sprite[3][40][53] = 1;cactus_sprite[3][40][54] = 1;cactus_sprite[3][40][55] = 1;cactus_sprite[3][40][56] = 1;cactus_sprite[3][40][57] = 1;cactus_sprite[3][40][58] = 1;cactus_sprite[3][40][59] = 1;cactus_sprite[3][40][60] = 1;cactus_sprite[3][40][61] = 1;cactus_sprite[3][40][62] = 1;cactus_sprite[3][40][63] = 1;cactus_sprite[3][41][28] = 1;cactus_sprite[3][41][29] = 1;cactus_sprite[3][41][30] = 1;cactus_sprite[3][41][31] = 1;cactus_sprite[3][41][32] = 1;cactus_sprite[3][41][33] = 1;cactus_sprite[3][41][34] = 1;cactus_sprite[3][41][35] = 1;cactus_sprite[3][41][36] = 1;cactus_sprite[3][41][37] = 1;cactus_sprite[3][41][38] = 1;cactus_sprite[3][41][39] = 1;cactus_sprite[3][41][40] = 1;cactus_sprite[3][41][41] = 1;cactus_sprite[3][41][42] = 1;cactus_sprite[3][41][43] = 1;cactus_sprite[3][41][44] = 1;cactus_sprite[3][41][45] = 1;cactus_sprite[3][41][46] = 1;cactus_sprite[3][41][47] = 1;cactus_sprite[3][41][48] = 1;cactus_sprite[3][41][49] = 1;cactus_sprite[3][41][50] = 1;cactus_sprite[3][41][51] = 1;cactus_sprite[3][41][52] = 1;cactus_sprite[3][41][53] = 1;cactus_sprite[3][41][54] = 1;cactus_sprite[3][41][55] = 1;cactus_sprite[3][41][56] = 1;cactus_sprite[3][41][57] = 1;cactus_sprite[3][41][58] = 1;cactus_sprite[3][41][59] = 1;cactus_sprite[3][41][60] = 1;cactus_sprite[3][41][61] = 1;cactus_sprite[3][41][62] = 1;cactus_sprite[3][41][63] = 1;cactus_sprite[3][42][28] = 1;cactus_sprite[3][42][29] = 1;cactus_sprite[3][42][30] = 1;cactus_sprite[3][42][31] = 1;cactus_sprite[3][42][32] = 1;cactus_sprite[3][42][33] = 1;cactus_sprite[3][42][34] = 1;cactus_sprite[3][42][35] = 1;cactus_sprite[3][42][36] = 1;cactus_sprite[3][42][37] = 1;cactus_sprite[3][42][38] = 1;cactus_sprite[3][42][39] = 1;cactus_sprite[3][42][40] = 1;cactus_sprite[3][42][41] = 1;cactus_sprite[3][42][42] = 1;cactus_sprite[3][42][43] = 1;cactus_sprite[3][42][44] = 1;cactus_sprite[3][42][45] = 1;cactus_sprite[3][42][46] = 1;cactus_sprite[3][42][47] = 1;cactus_sprite[3][42][48] = 1;cactus_sprite[3][42][49] = 1;cactus_sprite[3][42][50] = 1;cactus_sprite[3][42][51] = 1;cactus_sprite[3][42][52] = 1;cactus_sprite[3][42][53] = 1;cactus_sprite[3][42][54] = 1;cactus_sprite[3][42][55] = 1;cactus_sprite[3][42][56] = 1;cactus_sprite[3][42][57] = 1;cactus_sprite[3][42][58] = 1;cactus_sprite[3][42][59] = 1;cactus_sprite[3][42][60] = 1;cactus_sprite[3][42][61] = 1;cactus_sprite[3][43][28] = 1;cactus_sprite[3][43][29] = 1;cactus_sprite[3][43][30] = 1;cactus_sprite[3][43][31] = 1;cactus_sprite[3][43][32] = 1;cactus_sprite[3][43][33] = 1;cactus_sprite[3][43][34] = 1;cactus_sprite[3][43][35] = 1;cactus_sprite[3][43][36] = 1;cactus_sprite[3][43][37] = 1;cactus_sprite[3][43][38] = 1;cactus_sprite[3][43][39] = 1;cactus_sprite[3][43][40] = 1;cactus_sprite[3][43][41] = 1;cactus_sprite[3][43][42] = 1;cactus_sprite[3][43][43] = 1;cactus_sprite[3][43][44] = 1;cactus_sprite[3][43][45] = 1;cactus_sprite[3][43][46] = 1;cactus_sprite[3][43][47] = 1;cactus_sprite[3][43][48] = 1;cactus_sprite[3][43][49] = 1;cactus_sprite[3][43][50] = 1;cactus_sprite[3][43][51] = 1;cactus_sprite[3][43][52] = 1;cactus_sprite[3][43][53] = 1;cactus_sprite[3][43][54] = 1;cactus_sprite[3][43][55] = 1;cactus_sprite[3][43][56] = 1;cactus_sprite[3][43][57] = 1;cactus_sprite[3][43][58] = 1;cactus_sprite[3][43][59] = 1;cactus_sprite[3][43][60] = 1;cactus_sprite[3][43][61] = 1;cactus_sprite[3][44][30] = 1;cactus_sprite[3][44][31] = 1;cactus_sprite[3][44][32] = 1;cactus_sprite[3][44][33] = 1;cactus_sprite[3][44][34] = 1;cactus_sprite[3][44][35] = 1;cactus_sprite[3][44][36] = 1;cactus_sprite[3][44][37] = 1;cactus_sprite[3][44][38] = 1;cactus_sprite[3][44][39] = 1;cactus_sprite[3][44][40] = 1;cactus_sprite[3][44][41] = 1;cactus_sprite[3][44][42] = 1;cactus_sprite[3][44][43] = 1;cactus_sprite[3][44][44] = 1;cactus_sprite[3][44][45] = 1;cactus_sprite[3][44][46] = 1;cactus_sprite[3][44][47] = 1;cactus_sprite[3][44][48] = 1;cactus_sprite[3][44][49] = 1;cactus_sprite[3][44][50] = 1;cactus_sprite[3][44][51] = 1;cactus_sprite[3][44][52] = 1;cactus_sprite[3][44][53] = 1;cactus_sprite[3][44][54] = 1;cactus_sprite[3][44][55] = 1;cactus_sprite[3][44][56] = 1;cactus_sprite[3][44][57] = 1;cactus_sprite[3][44][58] = 1;cactus_sprite[3][44][59] = 1;cactus_sprite[3][45][30] = 1;cactus_sprite[3][45][31] = 1;cactus_sprite[3][45][32] = 1;cactus_sprite[3][45][33] = 1;cactus_sprite[3][45][34] = 1;cactus_sprite[3][45][35] = 1;cactus_sprite[3][45][36] = 1;cactus_sprite[3][45][37] = 1;cactus_sprite[3][45][38] = 1;cactus_sprite[3][45][39] = 1;cactus_sprite[3][45][40] = 1;cactus_sprite[3][45][41] = 1;cactus_sprite[3][45][42] = 1;cactus_sprite[3][45][43] = 1;cactus_sprite[3][45][44] = 1;cactus_sprite[3][45][45] = 1;cactus_sprite[3][45][46] = 1;cactus_sprite[3][45][47] = 1;cactus_sprite[3][45][48] = 1;cactus_sprite[3][45][49] = 1;cactus_sprite[3][45][50] = 1;cactus_sprite[3][45][51] = 1;cactus_sprite[3][45][52] = 1;cactus_sprite[3][45][53] = 1;cactus_sprite[3][45][54] = 1;cactus_sprite[3][45][55] = 1;cactus_sprite[3][45][56] = 1;cactus_sprite[3][45][57] = 1;cactus_sprite[3][45][58] = 1;cactus_sprite[3][45][59] = 1;
	cactus_sprite[4][2][41] = 1;cactus_sprite[4][2][42] = 1;cactus_sprite[4][2][43] = 1;cactus_sprite[4][2][44] = 1;cactus_sprite[4][2][45] = 1;cactus_sprite[4][2][46] = 1;cactus_sprite[4][2][47] = 1;cactus_sprite[4][2][48] = 1;cactus_sprite[4][2][49] = 1;cactus_sprite[4][2][50] = 1;cactus_sprite[4][2][51] = 1;cactus_sprite[4][2][52] = 1;cactus_sprite[4][2][53] = 1;cactus_sprite[4][2][54] = 1;cactus_sprite[4][2][55] = 1;cactus_sprite[4][2][56] = 1;cactus_sprite[4][2][57] = 1;cactus_sprite[4][2][58] = 1;cactus_sprite[4][2][59] = 1;cactus_sprite[4][2][60] = 1;cactus_sprite[4][2][61] = 1;cactus_sprite[4][2][62] = 1;cactus_sprite[4][2][63] = 1;cactus_sprite[4][2][64] = 1;cactus_sprite[4][2][65] = 1;cactus_sprite[4][2][66] = 1;cactus_sprite[4][3][41] = 1;cactus_sprite[4][3][42] = 1;cactus_sprite[4][3][43] = 1;cactus_sprite[4][3][44] = 1;cactus_sprite[4][3][45] = 1;cactus_sprite[4][3][46] = 1;cactus_sprite[4][3][47] = 1;cactus_sprite[4][3][48] = 1;cactus_sprite[4][3][49] = 1;cactus_sprite[4][3][50] = 1;cactus_sprite[4][3][51] = 1;cactus_sprite[4][3][52] = 1;cactus_sprite[4][3][53] = 1;cactus_sprite[4][3][54] = 1;cactus_sprite[4][3][55] = 1;cactus_sprite[4][3][56] = 1;cactus_sprite[4][3][57] = 1;cactus_sprite[4][3][58] = 1;cactus_sprite[4][3][59] = 1;cactus_sprite[4][3][60] = 1;cactus_sprite[4][3][61] = 1;cactus_sprite[4][3][62] = 1;cactus_sprite[4][3][63] = 1;cactus_sprite[4][3][64] = 1;cactus_sprite[4][3][65] = 1;cactus_sprite[4][3][66] = 1;cactus_sprite[4][4][39] = 1;cactus_sprite[4][4][40] = 1;cactus_sprite[4][4][41] = 1;cactus_sprite[4][4][42] = 1;cactus_sprite[4][4][43] = 1;cactus_sprite[4][4][44] = 1;cactus_sprite[4][4][45] = 1;cactus_sprite[4][4][46] = 1;cactus_sprite[4][4][47] = 1;cactus_sprite[4][4][48] = 1;cactus_sprite[4][4][49] = 1;cactus_sprite[4][4][50] = 1;cactus_sprite[4][4][51] = 1;cactus_sprite[4][4][52] = 1;cactus_sprite[4][4][53] = 1;cactus_sprite[4][4][54] = 1;cactus_sprite[4][4][55] = 1;cactus_sprite[4][4][56] = 1;cactus_sprite[4][4][57] = 1;cactus_sprite[4][4][58] = 1;cactus_sprite[4][4][59] = 1;cactus_sprite[4][4][60] = 1;cactus_sprite[4][4][61] = 1;cactus_sprite[4][4][62] = 1;cactus_sprite[4][4][63] = 1;cactus_sprite[4][4][64] = 1;cactus_sprite[4][4][65] = 1;cactus_sprite[4][4][66] = 1;cactus_sprite[4][4][67] = 1;cactus_sprite[4][4][68] = 1;cactus_sprite[4][5][39] = 1;cactus_sprite[4][5][40] = 1;cactus_sprite[4][5][41] = 1;cactus_sprite[4][5][42] = 1;cactus_sprite[4][5][43] = 1;cactus_sprite[4][5][44] = 1;cactus_sprite[4][5][45] = 1;cactus_sprite[4][5][46] = 1;cactus_sprite[4][5][47] = 1;cactus_sprite[4][5][48] = 1;cactus_sprite[4][5][49] = 1;cactus_sprite[4][5][50] = 1;cactus_sprite[4][5][51] = 1;cactus_sprite[4][5][52] = 1;cactus_sprite[4][5][53] = 1;cactus_sprite[4][5][54] = 1;cactus_sprite[4][5][55] = 1;cactus_sprite[4][5][56] = 1;cactus_sprite[4][5][57] = 1;cactus_sprite[4][5][58] = 1;cactus_sprite[4][5][59] = 1;cactus_sprite[4][5][60] = 1;cactus_sprite[4][5][61] = 1;cactus_sprite[4][5][62] = 1;cactus_sprite[4][5][63] = 1;cactus_sprite[4][5][64] = 1;cactus_sprite[4][5][65] = 1;cactus_sprite[4][5][66] = 1;cactus_sprite[4][5][67] = 1;cactus_sprite[4][5][68] = 1;cactus_sprite[4][6][39] = 1;cactus_sprite[4][6][40] = 1;cactus_sprite[4][6][41] = 1;cactus_sprite[4][6][42] = 1;cactus_sprite[4][6][43] = 1;cactus_sprite[4][6][44] = 1;cactus_sprite[4][6][45] = 1;cactus_sprite[4][6][46] = 1;cactus_sprite[4][6][47] = 1;cactus_sprite[4][6][48] = 1;cactus_sprite[4][6][49] = 1;cactus_sprite[4][6][50] = 1;cactus_sprite[4][6][51] = 1;cactus_sprite[4][6][52] = 1;cactus_sprite[4][6][53] = 1;cactus_sprite[4][6][54] = 1;cactus_sprite[4][6][55] = 1;cactus_sprite[4][6][56] = 1;cactus_sprite[4][6][57] = 1;cactus_sprite[4][6][58] = 1;cactus_sprite[4][6][59] = 1;cactus_sprite[4][6][60] = 1;cactus_sprite[4][6][61] = 1;cactus_sprite[4][6][62] = 1;cactus_sprite[4][6][63] = 1;cactus_sprite[4][6][64] = 1;cactus_sprite[4][6][65] = 1;cactus_sprite[4][6][66] = 1;cactus_sprite[4][6][67] = 1;cactus_sprite[4][6][68] = 1;cactus_sprite[4][6][69] = 1;cactus_sprite[4][6][70] = 1;cactus_sprite[4][7][39] = 1;cactus_sprite[4][7][40] = 1;cactus_sprite[4][7][41] = 1;cactus_sprite[4][7][42] = 1;cactus_sprite[4][7][43] = 1;cactus_sprite[4][7][44] = 1;cactus_sprite[4][7][45] = 1;cactus_sprite[4][7][46] = 1;cactus_sprite[4][7][47] = 1;cactus_sprite[4][7][48] = 1;cactus_sprite[4][7][49] = 1;cactus_sprite[4][7][50] = 1;cactus_sprite[4][7][51] = 1;cactus_sprite[4][7][52] = 1;cactus_sprite[4][7][53] = 1;cactus_sprite[4][7][54] = 1;cactus_sprite[4][7][55] = 1;cactus_sprite[4][7][56] = 1;cactus_sprite[4][7][57] = 1;cactus_sprite[4][7][58] = 1;cactus_sprite[4][7][59] = 1;cactus_sprite[4][7][60] = 1;cactus_sprite[4][7][61] = 1;cactus_sprite[4][7][62] = 1;cactus_sprite[4][7][63] = 1;cactus_sprite[4][7][64] = 1;cactus_sprite[4][7][65] = 1;cactus_sprite[4][7][66] = 1;cactus_sprite[4][7][67] = 1;cactus_sprite[4][7][68] = 1;cactus_sprite[4][7][69] = 1;cactus_sprite[4][7][70] = 1;cactus_sprite[4][8][41] = 1;cactus_sprite[4][8][42] = 1;cactus_sprite[4][8][43] = 1;cactus_sprite[4][8][44] = 1;cactus_sprite[4][8][45] = 1;cactus_sprite[4][8][46] = 1;cactus_sprite[4][8][47] = 1;cactus_sprite[4][8][48] = 1;cactus_sprite[4][8][49] = 1;cactus_sprite[4][8][50] = 1;cactus_sprite[4][8][51] = 1;cactus_sprite[4][8][52] = 1;cactus_sprite[4][8][53] = 1;cactus_sprite[4][8][54] = 1;cactus_sprite[4][8][55] = 1;cactus_sprite[4][8][56] = 1;cactus_sprite[4][8][57] = 1;cactus_sprite[4][8][58] = 1;cactus_sprite[4][8][59] = 1;cactus_sprite[4][8][60] = 1;cactus_sprite[4][8][61] = 1;cactus_sprite[4][8][62] = 1;cactus_sprite[4][8][63] = 1;cactus_sprite[4][8][64] = 1;cactus_sprite[4][8][65] = 1;cactus_sprite[4][8][66] = 1;cactus_sprite[4][8][67] = 1;cactus_sprite[4][8][68] = 1;cactus_sprite[4][8][69] = 1;cactus_sprite[4][8][70] = 1;cactus_sprite[4][8][71] = 1;cactus_sprite[4][8][72] = 1;cactus_sprite[4][9][41] = 1;cactus_sprite[4][9][42] = 1;cactus_sprite[4][9][43] = 1;cactus_sprite[4][9][44] = 1;cactus_sprite[4][9][45] = 1;cactus_sprite[4][9][46] = 1;cactus_sprite[4][9][47] = 1;cactus_sprite[4][9][48] = 1;cactus_sprite[4][9][49] = 1;cactus_sprite[4][9][50] = 1;cactus_sprite[4][9][51] = 1;cactus_sprite[4][9][52] = 1;cactus_sprite[4][9][53] = 1;cactus_sprite[4][9][54] = 1;cactus_sprite[4][9][55] = 1;cactus_sprite[4][9][56] = 1;cactus_sprite[4][9][57] = 1;cactus_sprite[4][9][58] = 1;cactus_sprite[4][9][59] = 1;cactus_sprite[4][9][60] = 1;cactus_sprite[4][9][61] = 1;cactus_sprite[4][9][62] = 1;cactus_sprite[4][9][63] = 1;cactus_sprite[4][9][64] = 1;cactus_sprite[4][9][65] = 1;cactus_sprite[4][9][66] = 1;cactus_sprite[4][9][67] = 1;cactus_sprite[4][9][68] = 1;cactus_sprite[4][9][69] = 1;cactus_sprite[4][9][70] = 1;cactus_sprite[4][9][71] = 1;cactus_sprite[4][9][72] = 1;cactus_sprite[4][10][65] = 1;cactus_sprite[4][10][66] = 1;cactus_sprite[4][10][67] = 1;cactus_sprite[4][10][68] = 1;cactus_sprite[4][10][69] = 1;cactus_sprite[4][10][70] = 1;cactus_sprite[4][10][71] = 1;cactus_sprite[4][10][72] = 1;cactus_sprite[4][11][65] = 1;cactus_sprite[4][11][66] = 1;cactus_sprite[4][11][67] = 1;cactus_sprite[4][11][68] = 1;cactus_sprite[4][11][69] = 1;cactus_sprite[4][11][70] = 1;cactus_sprite[4][11][71] = 1;cactus_sprite[4][11][72] = 1;cactus_sprite[4][12][65] = 1;cactus_sprite[4][12][66] = 1;cactus_sprite[4][12][67] = 1;cactus_sprite[4][12][68] = 1;cactus_sprite[4][12][69] = 1;cactus_sprite[4][12][70] = 1;cactus_sprite[4][12][71] = 1;cactus_sprite[4][12][72] = 1;cactus_sprite[4][13][65] = 1;cactus_sprite[4][13][66] = 1;cactus_sprite[4][13][67] = 1;cactus_sprite[4][13][68] = 1;cactus_sprite[4][13][69] = 1;cactus_sprite[4][13][70] = 1;cactus_sprite[4][13][71] = 1;cactus_sprite[4][13][72] = 1;cactus_sprite[4][14][13] = 1;cactus_sprite[4][14][14] = 1;cactus_sprite[4][14][15] = 1;cactus_sprite[4][14][16] = 1;cactus_sprite[4][14][17] = 1;cactus_sprite[4][14][18] = 1;cactus_sprite[4][14][19] = 1;cactus_sprite[4][14][20] = 1;cactus_sprite[4][14][21] = 1;cactus_sprite[4][14][22] = 1;cactus_sprite[4][14][23] = 1;cactus_sprite[4][14][24] = 1;cactus_sprite[4][14][25] = 1;cactus_sprite[4][14][26] = 1;cactus_sprite[4][14][27] = 1;cactus_sprite[4][14][28] = 1;cactus_sprite[4][14][29] = 1;cactus_sprite[4][14][30] = 1;cactus_sprite[4][14][31] = 1;cactus_sprite[4][14][32] = 1;cactus_sprite[4][14][33] = 1;cactus_sprite[4][14][34] = 1;cactus_sprite[4][14][35] = 1;cactus_sprite[4][14][36] = 1;cactus_sprite[4][14][37] = 1;cactus_sprite[4][14][38] = 1;cactus_sprite[4][14][39] = 1;cactus_sprite[4][14][40] = 1;cactus_sprite[4][14][41] = 1;cactus_sprite[4][14][42] = 1;cactus_sprite[4][14][43] = 1;cactus_sprite[4][14][44] = 1;cactus_sprite[4][14][45] = 1;cactus_sprite[4][14][46] = 1;cactus_sprite[4][14][47] = 1;cactus_sprite[4][14][48] = 1;cactus_sprite[4][14][49] = 1;cactus_sprite[4][14][50] = 1;cactus_sprite[4][14][51] = 1;cactus_sprite[4][14][52] = 1;cactus_sprite[4][14][53] = 1;cactus_sprite[4][14][54] = 1;cactus_sprite[4][14][55] = 1;cactus_sprite[4][14][56] = 1;cactus_sprite[4][14][57] = 1;cactus_sprite[4][14][58] = 1;cactus_sprite[4][14][59] = 1;cactus_sprite[4][14][60] = 1;cactus_sprite[4][14][61] = 1;cactus_sprite[4][14][62] = 1;cactus_sprite[4][14][63] = 1;cactus_sprite[4][14][64] = 1;cactus_sprite[4][14][65] = 1;cactus_sprite[4][14][66] = 1;cactus_sprite[4][14][67] = 1;cactus_sprite[4][14][68] = 1;cactus_sprite[4][14][69] = 1;cactus_sprite[4][14][70] = 1;cactus_sprite[4][14][71] = 1;cactus_sprite[4][14][72] = 1;cactus_sprite[4][14][73] = 1;cactus_sprite[4][14][74] = 1;cactus_sprite[4][14][75] = 1;cactus_sprite[4][14][76] = 1;cactus_sprite[4][14][77] = 1;cactus_sprite[4][14][78] = 1;cactus_sprite[4][14][79] = 1;cactus_sprite[4][14][80] = 1;cactus_sprite[4][14][81] = 1;cactus_sprite[4][14][82] = 1;cactus_sprite[4][14][83] = 1;cactus_sprite[4][14][84] = 1;cactus_sprite[4][14][85] = 1;cactus_sprite[4][14][86] = 1;cactus_sprite[4][14][87] = 1;cactus_sprite[4][14][88] = 1;cactus_sprite[4][14][89] = 1;cactus_sprite[4][14][90] = 1;cactus_sprite[4][14][91] = 1;cactus_sprite[4][14][92] = 1;cactus_sprite[4][14][93] = 1;cactus_sprite[4][14][94] = 1;cactus_sprite[4][14][95] = 1;cactus_sprite[4][14][96] = 1;cactus_sprite[4][14][97] = 1;cactus_sprite[4][14][98] = 1;cactus_sprite[4][14][99] = 1;cactus_sprite[4][15][13] = 1;cactus_sprite[4][15][14] = 1;cactus_sprite[4][15][15] = 1;cactus_sprite[4][15][16] = 1;cactus_sprite[4][15][17] = 1;cactus_sprite[4][15][18] = 1;cactus_sprite[4][15][19] = 1;cactus_sprite[4][15][20] = 1;cactus_sprite[4][15][21] = 1;cactus_sprite[4][15][22] = 1;cactus_sprite[4][15][23] = 1;cactus_sprite[4][15][24] = 1;cactus_sprite[4][15][25] = 1;cactus_sprite[4][15][26] = 1;cactus_sprite[4][15][27] = 1;cactus_sprite[4][15][28] = 1;cactus_sprite[4][15][29] = 1;cactus_sprite[4][15][30] = 1;cactus_sprite[4][15][31] = 1;cactus_sprite[4][15][32] = 1;cactus_sprite[4][15][33] = 1;cactus_sprite[4][15][34] = 1;cactus_sprite[4][15][35] = 1;cactus_sprite[4][15][36] = 1;cactus_sprite[4][15][37] = 1;cactus_sprite[4][15][38] = 1;cactus_sprite[4][15][39] = 1;cactus_sprite[4][15][40] = 1;cactus_sprite[4][15][41] = 1;cactus_sprite[4][15][42] = 1;cactus_sprite[4][15][43] = 1;cactus_sprite[4][15][44] = 1;cactus_sprite[4][15][45] = 1;cactus_sprite[4][15][46] = 1;cactus_sprite[4][15][47] = 1;cactus_sprite[4][15][48] = 1;cactus_sprite[4][15][49] = 1;cactus_sprite[4][15][50] = 1;cactus_sprite[4][15][51] = 1;cactus_sprite[4][15][52] = 1;cactus_sprite[4][15][53] = 1;cactus_sprite[4][15][54] = 1;cactus_sprite[4][15][55] = 1;cactus_sprite[4][15][56] = 1;cactus_sprite[4][15][57] = 1;cactus_sprite[4][15][58] = 1;cactus_sprite[4][15][59] = 1;cactus_sprite[4][15][60] = 1;cactus_sprite[4][15][61] = 1;cactus_sprite[4][15][62] = 1;cactus_sprite[4][15][63] = 1;cactus_sprite[4][15][64] = 1;cactus_sprite[4][15][65] = 1;cactus_sprite[4][15][66] = 1;cactus_sprite[4][15][67] = 1;cactus_sprite[4][15][68] = 1;cactus_sprite[4][15][69] = 1;cactus_sprite[4][15][70] = 1;cactus_sprite[4][15][71] = 1;cactus_sprite[4][15][72] = 1;cactus_sprite[4][15][73] = 1;cactus_sprite[4][15][74] = 1;cactus_sprite[4][15][75] = 1;cactus_sprite[4][15][76] = 1;cactus_sprite[4][15][77] = 1;cactus_sprite[4][15][78] = 1;cactus_sprite[4][15][79] = 1;cactus_sprite[4][15][80] = 1;cactus_sprite[4][15][81] = 1;cactus_sprite[4][15][82] = 1;cactus_sprite[4][15][83] = 1;cactus_sprite[4][15][84] = 1;cactus_sprite[4][15][85] = 1;cactus_sprite[4][15][86] = 1;cactus_sprite[4][15][87] = 1;cactus_sprite[4][15][88] = 1;cactus_sprite[4][15][89] = 1;cactus_sprite[4][15][90] = 1;cactus_sprite[4][15][91] = 1;cactus_sprite[4][15][92] = 1;cactus_sprite[4][15][93] = 1;cactus_sprite[4][15][94] = 1;cactus_sprite[4][15][95] = 1;cactus_sprite[4][15][96] = 1;cactus_sprite[4][15][97] = 1;cactus_sprite[4][15][98] = 1;cactus_sprite[4][15][99] = 1;cactus_sprite[4][16][11] = 1;cactus_sprite[4][16][12] = 1;cactus_sprite[4][16][13] = 1;cactus_sprite[4][16][14] = 1;cactus_sprite[4][16][15] = 1;cactus_sprite[4][16][16] = 1;cactus_sprite[4][16][17] = 1;cactus_sprite[4][16][18] = 1;cactus_sprite[4][16][19] = 1;cactus_sprite[4][16][20] = 1;cactus_sprite[4][16][21] = 1;cactus_sprite[4][16][22] = 1;cactus_sprite[4][16][23] = 1;cactus_sprite[4][16][24] = 1;cactus_sprite[4][16][25] = 1;cactus_sprite[4][16][26] = 1;cactus_sprite[4][16][27] = 1;cactus_sprite[4][16][28] = 1;cactus_sprite[4][16][29] = 1;cactus_sprite[4][16][30] = 1;cactus_sprite[4][16][31] = 1;cactus_sprite[4][16][32] = 1;cactus_sprite[4][16][33] = 1;cactus_sprite[4][16][34] = 1;cactus_sprite[4][16][35] = 1;cactus_sprite[4][16][36] = 1;cactus_sprite[4][16][37] = 1;cactus_sprite[4][16][38] = 1;cactus_sprite[4][16][39] = 1;cactus_sprite[4][16][40] = 1;cactus_sprite[4][16][41] = 1;cactus_sprite[4][16][42] = 1;cactus_sprite[4][16][43] = 1;cactus_sprite[4][16][44] = 1;cactus_sprite[4][16][45] = 1;cactus_sprite[4][16][46] = 1;cactus_sprite[4][16][47] = 1;cactus_sprite[4][16][48] = 1;cactus_sprite[4][16][49] = 1;cactus_sprite[4][16][50] = 1;cactus_sprite[4][16][51] = 1;cactus_sprite[4][16][52] = 1;cactus_sprite[4][16][53] = 1;cactus_sprite[4][16][54] = 1;cactus_sprite[4][16][55] = 1;cactus_sprite[4][16][56] = 1;cactus_sprite[4][16][57] = 1;cactus_sprite[4][16][58] = 1;cactus_sprite[4][16][59] = 1;cactus_sprite[4][16][60] = 1;cactus_sprite[4][16][61] = 1;cactus_sprite[4][16][62] = 1;cactus_sprite[4][16][63] = 1;cactus_sprite[4][16][64] = 1;cactus_sprite[4][16][65] = 1;cactus_sprite[4][16][66] = 1;cactus_sprite[4][16][67] = 1;cactus_sprite[4][16][68] = 1;cactus_sprite[4][16][69] = 1;cactus_sprite[4][16][70] = 1;cactus_sprite[4][16][71] = 1;cactus_sprite[4][16][72] = 1;cactus_sprite[4][16][73] = 1;cactus_sprite[4][16][74] = 1;cactus_sprite[4][16][75] = 1;cactus_sprite[4][16][76] = 1;cactus_sprite[4][16][77] = 1;cactus_sprite[4][16][78] = 1;cactus_sprite[4][16][79] = 1;cactus_sprite[4][16][80] = 1;cactus_sprite[4][16][81] = 1;cactus_sprite[4][16][82] = 1;cactus_sprite[4][16][83] = 1;cactus_sprite[4][16][84] = 1;cactus_sprite[4][16][85] = 1;cactus_sprite[4][16][86] = 1;cactus_sprite[4][16][87] = 1;cactus_sprite[4][16][88] = 1;cactus_sprite[4][16][89] = 1;cactus_sprite[4][16][90] = 1;cactus_sprite[4][16][91] = 1;cactus_sprite[4][16][92] = 1;cactus_sprite[4][16][93] = 1;cactus_sprite[4][16][94] = 1;cactus_sprite[4][16][95] = 1;cactus_sprite[4][16][96] = 1;cactus_sprite[4][16][97] = 1;cactus_sprite[4][16][98] = 1;cactus_sprite[4][16][99] = 1;cactus_sprite[4][17][11] = 1;cactus_sprite[4][17][12] = 1;cactus_sprite[4][17][13] = 1;cactus_sprite[4][17][14] = 1;cactus_sprite[4][17][15] = 1;cactus_sprite[4][17][16] = 1;cactus_sprite[4][17][17] = 1;cactus_sprite[4][17][18] = 1;cactus_sprite[4][17][19] = 1;cactus_sprite[4][17][20] = 1;cactus_sprite[4][17][21] = 1;cactus_sprite[4][17][22] = 1;cactus_sprite[4][17][23] = 1;cactus_sprite[4][17][24] = 1;cactus_sprite[4][17][25] = 1;cactus_sprite[4][17][26] = 1;cactus_sprite[4][17][27] = 1;cactus_sprite[4][17][28] = 1;cactus_sprite[4][17][29] = 1;cactus_sprite[4][17][30] = 1;cactus_sprite[4][17][31] = 1;cactus_sprite[4][17][32] = 1;cactus_sprite[4][17][33] = 1;cactus_sprite[4][17][34] = 1;cactus_sprite[4][17][35] = 1;cactus_sprite[4][17][36] = 1;cactus_sprite[4][17][37] = 1;cactus_sprite[4][17][38] = 1;cactus_sprite[4][17][39] = 1;cactus_sprite[4][17][40] = 1;cactus_sprite[4][17][41] = 1;cactus_sprite[4][17][42] = 1;cactus_sprite[4][17][43] = 1;cactus_sprite[4][17][44] = 1;cactus_sprite[4][17][45] = 1;cactus_sprite[4][17][46] = 1;cactus_sprite[4][17][47] = 1;cactus_sprite[4][17][48] = 1;cactus_sprite[4][17][49] = 1;cactus_sprite[4][17][50] = 1;cactus_sprite[4][17][51] = 1;cactus_sprite[4][17][52] = 1;cactus_sprite[4][17][53] = 1;cactus_sprite[4][17][54] = 1;cactus_sprite[4][17][55] = 1;cactus_sprite[4][17][56] = 1;cactus_sprite[4][17][57] = 1;cactus_sprite[4][17][58] = 1;cactus_sprite[4][17][59] = 1;cactus_sprite[4][17][60] = 1;cactus_sprite[4][17][61] = 1;cactus_sprite[4][17][62] = 1;cactus_sprite[4][17][63] = 1;cactus_sprite[4][17][64] = 1;cactus_sprite[4][17][65] = 1;cactus_sprite[4][17][66] = 1;cactus_sprite[4][17][67] = 1;cactus_sprite[4][17][68] = 1;cactus_sprite[4][17][69] = 1;cactus_sprite[4][17][70] = 1;cactus_sprite[4][17][71] = 1;cactus_sprite[4][17][72] = 1;cactus_sprite[4][17][73] = 1;cactus_sprite[4][17][74] = 1;cactus_sprite[4][17][75] = 1;cactus_sprite[4][17][76] = 1;cactus_sprite[4][17][77] = 1;cactus_sprite[4][17][78] = 1;cactus_sprite[4][17][79] = 1;cactus_sprite[4][17][80] = 1;cactus_sprite[4][17][81] = 1;cactus_sprite[4][17][82] = 1;cactus_sprite[4][17][83] = 1;cactus_sprite[4][17][84] = 1;cactus_sprite[4][17][85] = 1;cactus_sprite[4][17][86] = 1;cactus_sprite[4][17][87] = 1;cactus_sprite[4][17][88] = 1;cactus_sprite[4][17][89] = 1;cactus_sprite[4][17][90] = 1;cactus_sprite[4][17][91] = 1;cactus_sprite[4][17][92] = 1;cactus_sprite[4][17][93] = 1;cactus_sprite[4][17][94] = 1;cactus_sprite[4][17][95] = 1;cactus_sprite[4][17][96] = 1;cactus_sprite[4][17][97] = 1;cactus_sprite[4][17][98] = 1;cactus_sprite[4][17][99] = 1;cactus_sprite[4][18][11] = 1;cactus_sprite[4][18][12] = 1;cactus_sprite[4][18][13] = 1;cactus_sprite[4][18][14] = 1;cactus_sprite[4][18][15] = 1;cactus_sprite[4][18][16] = 1;cactus_sprite[4][18][17] = 1;cactus_sprite[4][18][18] = 1;cactus_sprite[4][18][19] = 1;cactus_sprite[4][18][20] = 1;cactus_sprite[4][18][21] = 1;cactus_sprite[4][18][22] = 1;cactus_sprite[4][18][23] = 1;cactus_sprite[4][18][24] = 1;cactus_sprite[4][18][25] = 1;cactus_sprite[4][18][26] = 1;cactus_sprite[4][18][27] = 1;cactus_sprite[4][18][28] = 1;cactus_sprite[4][18][29] = 1;cactus_sprite[4][18][30] = 1;cactus_sprite[4][18][31] = 1;cactus_sprite[4][18][32] = 1;cactus_sprite[4][18][33] = 1;cactus_sprite[4][18][34] = 1;cactus_sprite[4][18][35] = 1;cactus_sprite[4][18][36] = 1;cactus_sprite[4][18][37] = 1;cactus_sprite[4][18][38] = 1;cactus_sprite[4][18][39] = 1;cactus_sprite[4][18][40] = 1;cactus_sprite[4][18][41] = 1;cactus_sprite[4][18][42] = 1;cactus_sprite[4][18][43] = 1;cactus_sprite[4][18][44] = 1;cactus_sprite[4][18][45] = 1;cactus_sprite[4][18][46] = 1;cactus_sprite[4][18][47] = 1;cactus_sprite[4][18][48] = 1;cactus_sprite[4][18][49] = 1;cactus_sprite[4][18][50] = 1;cactus_sprite[4][18][51] = 1;cactus_sprite[4][18][52] = 1;cactus_sprite[4][18][53] = 1;cactus_sprite[4][18][54] = 1;cactus_sprite[4][18][55] = 1;cactus_sprite[4][18][56] = 1;cactus_sprite[4][18][57] = 1;cactus_sprite[4][18][58] = 1;cactus_sprite[4][18][59] = 1;cactus_sprite[4][18][60] = 1;cactus_sprite[4][18][61] = 1;cactus_sprite[4][18][62] = 1;cactus_sprite[4][18][63] = 1;cactus_sprite[4][18][64] = 1;cactus_sprite[4][18][65] = 1;cactus_sprite[4][18][66] = 1;cactus_sprite[4][18][67] = 1;cactus_sprite[4][18][68] = 1;cactus_sprite[4][18][69] = 1;cactus_sprite[4][18][70] = 1;cactus_sprite[4][18][71] = 1;cactus_sprite[4][18][72] = 1;cactus_sprite[4][18][73] = 1;cactus_sprite[4][18][74] = 1;cactus_sprite[4][18][75] = 1;cactus_sprite[4][18][76] = 1;cactus_sprite[4][18][77] = 1;cactus_sprite[4][18][78] = 1;cactus_sprite[4][18][79] = 1;cactus_sprite[4][18][80] = 1;cactus_sprite[4][18][81] = 1;cactus_sprite[4][18][82] = 1;cactus_sprite[4][18][83] = 1;cactus_sprite[4][18][84] = 1;cactus_sprite[4][18][85] = 1;cactus_sprite[4][18][86] = 1;cactus_sprite[4][18][87] = 1;cactus_sprite[4][18][88] = 1;cactus_sprite[4][18][89] = 1;cactus_sprite[4][18][90] = 1;cactus_sprite[4][18][91] = 1;cactus_sprite[4][18][92] = 1;cactus_sprite[4][18][93] = 1;cactus_sprite[4][18][94] = 1;cactus_sprite[4][18][95] = 1;cactus_sprite[4][18][96] = 1;cactus_sprite[4][18][97] = 1;cactus_sprite[4][18][98] = 1;cactus_sprite[4][18][99] = 1;cactus_sprite[4][19][11] = 1;cactus_sprite[4][19][12] = 1;cactus_sprite[4][19][13] = 1;cactus_sprite[4][19][14] = 1;cactus_sprite[4][19][15] = 1;cactus_sprite[4][19][16] = 1;cactus_sprite[4][19][17] = 1;cactus_sprite[4][19][18] = 1;cactus_sprite[4][19][19] = 1;cactus_sprite[4][19][20] = 1;cactus_sprite[4][19][21] = 1;cactus_sprite[4][19][22] = 1;cactus_sprite[4][19][23] = 1;cactus_sprite[4][19][24] = 1;cactus_sprite[4][19][25] = 1;cactus_sprite[4][19][26] = 1;cactus_sprite[4][19][27] = 1;cactus_sprite[4][19][28] = 1;cactus_sprite[4][19][29] = 1;cactus_sprite[4][19][30] = 1;cactus_sprite[4][19][31] = 1;cactus_sprite[4][19][32] = 1;cactus_sprite[4][19][33] = 1;cactus_sprite[4][19][34] = 1;cactus_sprite[4][19][35] = 1;cactus_sprite[4][19][36] = 1;cactus_sprite[4][19][37] = 1;cactus_sprite[4][19][38] = 1;cactus_sprite[4][19][39] = 1;cactus_sprite[4][19][40] = 1;cactus_sprite[4][19][41] = 1;cactus_sprite[4][19][42] = 1;cactus_sprite[4][19][43] = 1;cactus_sprite[4][19][44] = 1;cactus_sprite[4][19][45] = 1;cactus_sprite[4][19][46] = 1;cactus_sprite[4][19][47] = 1;cactus_sprite[4][19][48] = 1;cactus_sprite[4][19][49] = 1;cactus_sprite[4][19][50] = 1;cactus_sprite[4][19][51] = 1;cactus_sprite[4][19][52] = 1;cactus_sprite[4][19][53] = 1;cactus_sprite[4][19][54] = 1;cactus_sprite[4][19][55] = 1;cactus_sprite[4][19][56] = 1;cactus_sprite[4][19][57] = 1;cactus_sprite[4][19][58] = 1;cactus_sprite[4][19][59] = 1;cactus_sprite[4][19][60] = 1;cactus_sprite[4][19][61] = 1;cactus_sprite[4][19][62] = 1;cactus_sprite[4][19][63] = 1;cactus_sprite[4][19][64] = 1;cactus_sprite[4][19][65] = 1;cactus_sprite[4][19][66] = 1;cactus_sprite[4][19][67] = 1;cactus_sprite[4][19][68] = 1;cactus_sprite[4][19][69] = 1;cactus_sprite[4][19][70] = 1;cactus_sprite[4][19][71] = 1;cactus_sprite[4][19][72] = 1;cactus_sprite[4][19][73] = 1;cactus_sprite[4][19][74] = 1;cactus_sprite[4][19][75] = 1;cactus_sprite[4][19][76] = 1;cactus_sprite[4][19][77] = 1;cactus_sprite[4][19][78] = 1;cactus_sprite[4][19][79] = 1;cactus_sprite[4][19][80] = 1;cactus_sprite[4][19][81] = 1;cactus_sprite[4][19][82] = 1;cactus_sprite[4][19][83] = 1;cactus_sprite[4][19][84] = 1;cactus_sprite[4][19][85] = 1;cactus_sprite[4][19][86] = 1;cactus_sprite[4][19][87] = 1;cactus_sprite[4][19][88] = 1;cactus_sprite[4][19][89] = 1;cactus_sprite[4][19][90] = 1;cactus_sprite[4][19][91] = 1;cactus_sprite[4][19][92] = 1;cactus_sprite[4][19][93] = 1;cactus_sprite[4][19][94] = 1;cactus_sprite[4][19][95] = 1;cactus_sprite[4][19][96] = 1;cactus_sprite[4][19][97] = 1;cactus_sprite[4][19][98] = 1;cactus_sprite[4][19][99] = 1;cactus_sprite[4][20][11] = 1;cactus_sprite[4][20][12] = 1;cactus_sprite[4][20][13] = 1;cactus_sprite[4][20][14] = 1;cactus_sprite[4][20][15] = 1;cactus_sprite[4][20][16] = 1;cactus_sprite[4][20][17] = 1;cactus_sprite[4][20][18] = 1;cactus_sprite[4][20][19] = 1;cactus_sprite[4][20][20] = 1;cactus_sprite[4][20][21] = 1;cactus_sprite[4][20][22] = 1;cactus_sprite[4][20][23] = 1;cactus_sprite[4][20][24] = 1;cactus_sprite[4][20][25] = 1;cactus_sprite[4][20][26] = 1;cactus_sprite[4][20][27] = 1;cactus_sprite[4][20][28] = 1;cactus_sprite[4][20][29] = 1;cactus_sprite[4][20][30] = 1;cactus_sprite[4][20][31] = 1;cactus_sprite[4][20][32] = 1;cactus_sprite[4][20][33] = 1;cactus_sprite[4][20][34] = 1;cactus_sprite[4][20][35] = 1;cactus_sprite[4][20][36] = 1;cactus_sprite[4][20][37] = 1;cactus_sprite[4][20][38] = 1;cactus_sprite[4][20][39] = 1;cactus_sprite[4][20][40] = 1;cactus_sprite[4][20][41] = 1;cactus_sprite[4][20][42] = 1;cactus_sprite[4][20][43] = 1;cactus_sprite[4][20][44] = 1;cactus_sprite[4][20][45] = 1;cactus_sprite[4][20][46] = 1;cactus_sprite[4][20][47] = 1;cactus_sprite[4][20][48] = 1;cactus_sprite[4][20][49] = 1;cactus_sprite[4][20][50] = 1;cactus_sprite[4][20][51] = 1;cactus_sprite[4][20][52] = 1;cactus_sprite[4][20][53] = 1;cactus_sprite[4][20][54] = 1;cactus_sprite[4][20][55] = 1;cactus_sprite[4][20][56] = 1;cactus_sprite[4][20][57] = 1;cactus_sprite[4][20][58] = 1;cactus_sprite[4][20][59] = 1;cactus_sprite[4][20][60] = 1;cactus_sprite[4][20][61] = 1;cactus_sprite[4][20][62] = 1;cactus_sprite[4][20][63] = 1;cactus_sprite[4][20][64] = 1;cactus_sprite[4][20][65] = 1;cactus_sprite[4][20][66] = 1;cactus_sprite[4][20][67] = 1;cactus_sprite[4][20][68] = 1;cactus_sprite[4][20][69] = 1;cactus_sprite[4][20][70] = 1;cactus_sprite[4][20][71] = 1;cactus_sprite[4][20][72] = 1;cactus_sprite[4][20][73] = 1;cactus_sprite[4][20][74] = 1;cactus_sprite[4][20][75] = 1;cactus_sprite[4][20][76] = 1;cactus_sprite[4][20][77] = 1;cactus_sprite[4][20][78] = 1;cactus_sprite[4][20][79] = 1;cactus_sprite[4][20][80] = 1;cactus_sprite[4][20][81] = 1;cactus_sprite[4][20][82] = 1;cactus_sprite[4][20][83] = 1;cactus_sprite[4][20][84] = 1;cactus_sprite[4][20][85] = 1;cactus_sprite[4][20][86] = 1;cactus_sprite[4][20][87] = 1;cactus_sprite[4][20][88] = 1;cactus_sprite[4][20][89] = 1;cactus_sprite[4][20][90] = 1;cactus_sprite[4][20][91] = 1;cactus_sprite[4][20][92] = 1;cactus_sprite[4][20][93] = 1;cactus_sprite[4][20][94] = 1;cactus_sprite[4][20][95] = 1;cactus_sprite[4][20][96] = 1;cactus_sprite[4][20][97] = 1;cactus_sprite[4][20][98] = 1;cactus_sprite[4][20][99] = 1;cactus_sprite[4][21][11] = 1;cactus_sprite[4][21][12] = 1;cactus_sprite[4][21][13] = 1;cactus_sprite[4][21][14] = 1;cactus_sprite[4][21][15] = 1;cactus_sprite[4][21][16] = 1;cactus_sprite[4][21][17] = 1;cactus_sprite[4][21][18] = 1;cactus_sprite[4][21][19] = 1;cactus_sprite[4][21][20] = 1;cactus_sprite[4][21][21] = 1;cactus_sprite[4][21][22] = 1;cactus_sprite[4][21][23] = 1;cactus_sprite[4][21][24] = 1;cactus_sprite[4][21][25] = 1;cactus_sprite[4][21][26] = 1;cactus_sprite[4][21][27] = 1;cactus_sprite[4][21][28] = 1;cactus_sprite[4][21][29] = 1;cactus_sprite[4][21][30] = 1;cactus_sprite[4][21][31] = 1;cactus_sprite[4][21][32] = 1;cactus_sprite[4][21][33] = 1;cactus_sprite[4][21][34] = 1;cactus_sprite[4][21][35] = 1;cactus_sprite[4][21][36] = 1;cactus_sprite[4][21][37] = 1;cactus_sprite[4][21][38] = 1;cactus_sprite[4][21][39] = 1;cactus_sprite[4][21][40] = 1;cactus_sprite[4][21][41] = 1;cactus_sprite[4][21][42] = 1;cactus_sprite[4][21][43] = 1;cactus_sprite[4][21][44] = 1;cactus_sprite[4][21][45] = 1;cactus_sprite[4][21][46] = 1;cactus_sprite[4][21][47] = 1;cactus_sprite[4][21][48] = 1;cactus_sprite[4][21][49] = 1;cactus_sprite[4][21][50] = 1;cactus_sprite[4][21][51] = 1;cactus_sprite[4][21][52] = 1;cactus_sprite[4][21][53] = 1;cactus_sprite[4][21][54] = 1;cactus_sprite[4][21][55] = 1;cactus_sprite[4][21][56] = 1;cactus_sprite[4][21][57] = 1;cactus_sprite[4][21][58] = 1;cactus_sprite[4][21][59] = 1;cactus_sprite[4][21][60] = 1;cactus_sprite[4][21][61] = 1;cactus_sprite[4][21][62] = 1;cactus_sprite[4][21][63] = 1;cactus_sprite[4][21][64] = 1;cactus_sprite[4][21][65] = 1;cactus_sprite[4][21][66] = 1;cactus_sprite[4][21][67] = 1;cactus_sprite[4][21][68] = 1;cactus_sprite[4][21][69] = 1;cactus_sprite[4][21][70] = 1;cactus_sprite[4][21][71] = 1;cactus_sprite[4][21][72] = 1;cactus_sprite[4][21][73] = 1;cactus_sprite[4][21][74] = 1;cactus_sprite[4][21][75] = 1;cactus_sprite[4][21][76] = 1;cactus_sprite[4][21][77] = 1;cactus_sprite[4][21][78] = 1;cactus_sprite[4][21][79] = 1;cactus_sprite[4][21][80] = 1;cactus_sprite[4][21][81] = 1;cactus_sprite[4][21][82] = 1;cactus_sprite[4][21][83] = 1;cactus_sprite[4][21][84] = 1;cactus_sprite[4][21][85] = 1;cactus_sprite[4][21][86] = 1;cactus_sprite[4][21][87] = 1;cactus_sprite[4][21][88] = 1;cactus_sprite[4][21][89] = 1;cactus_sprite[4][21][90] = 1;cactus_sprite[4][21][91] = 1;cactus_sprite[4][21][92] = 1;cactus_sprite[4][21][93] = 1;cactus_sprite[4][21][94] = 1;cactus_sprite[4][21][95] = 1;cactus_sprite[4][21][96] = 1;cactus_sprite[4][21][97] = 1;cactus_sprite[4][21][98] = 1;cactus_sprite[4][21][99] = 1;cactus_sprite[4][22][13] = 1;cactus_sprite[4][22][14] = 1;cactus_sprite[4][22][15] = 1;cactus_sprite[4][22][16] = 1;cactus_sprite[4][22][17] = 1;cactus_sprite[4][22][18] = 1;cactus_sprite[4][22][19] = 1;cactus_sprite[4][22][20] = 1;cactus_sprite[4][22][21] = 1;cactus_sprite[4][22][22] = 1;cactus_sprite[4][22][23] = 1;cactus_sprite[4][22][24] = 1;cactus_sprite[4][22][25] = 1;cactus_sprite[4][22][26] = 1;cactus_sprite[4][22][27] = 1;cactus_sprite[4][22][28] = 1;cactus_sprite[4][22][29] = 1;cactus_sprite[4][22][30] = 1;cactus_sprite[4][22][31] = 1;cactus_sprite[4][22][32] = 1;cactus_sprite[4][22][33] = 1;cactus_sprite[4][22][34] = 1;cactus_sprite[4][22][35] = 1;cactus_sprite[4][22][36] = 1;cactus_sprite[4][22][37] = 1;cactus_sprite[4][22][38] = 1;cactus_sprite[4][22][39] = 1;cactus_sprite[4][22][40] = 1;cactus_sprite[4][22][41] = 1;cactus_sprite[4][22][42] = 1;cactus_sprite[4][22][43] = 1;cactus_sprite[4][22][44] = 1;cactus_sprite[4][22][45] = 1;cactus_sprite[4][22][46] = 1;cactus_sprite[4][22][47] = 1;cactus_sprite[4][22][48] = 1;cactus_sprite[4][22][49] = 1;cactus_sprite[4][22][50] = 1;cactus_sprite[4][22][51] = 1;cactus_sprite[4][22][52] = 1;cactus_sprite[4][22][53] = 1;cactus_sprite[4][22][54] = 1;cactus_sprite[4][22][55] = 1;cactus_sprite[4][22][56] = 1;cactus_sprite[4][22][57] = 1;cactus_sprite[4][22][58] = 1;cactus_sprite[4][22][59] = 1;cactus_sprite[4][22][60] = 1;cactus_sprite[4][22][61] = 1;cactus_sprite[4][22][62] = 1;cactus_sprite[4][22][63] = 1;cactus_sprite[4][22][64] = 1;cactus_sprite[4][22][65] = 1;cactus_sprite[4][22][66] = 1;cactus_sprite[4][22][67] = 1;cactus_sprite[4][22][68] = 1;cactus_sprite[4][22][69] = 1;cactus_sprite[4][22][70] = 1;cactus_sprite[4][22][71] = 1;cactus_sprite[4][22][72] = 1;cactus_sprite[4][22][73] = 1;cactus_sprite[4][22][74] = 1;cactus_sprite[4][22][75] = 1;cactus_sprite[4][22][76] = 1;cactus_sprite[4][22][77] = 1;cactus_sprite[4][22][78] = 1;cactus_sprite[4][22][79] = 1;cactus_sprite[4][22][80] = 1;cactus_sprite[4][22][81] = 1;cactus_sprite[4][22][82] = 1;cactus_sprite[4][22][83] = 1;cactus_sprite[4][22][84] = 1;cactus_sprite[4][22][85] = 1;cactus_sprite[4][22][86] = 1;cactus_sprite[4][22][87] = 1;cactus_sprite[4][22][88] = 1;cactus_sprite[4][22][89] = 1;cactus_sprite[4][22][90] = 1;cactus_sprite[4][22][91] = 1;cactus_sprite[4][22][92] = 1;cactus_sprite[4][22][93] = 1;cactus_sprite[4][22][94] = 1;cactus_sprite[4][22][95] = 1;cactus_sprite[4][22][96] = 1;cactus_sprite[4][22][97] = 1;cactus_sprite[4][22][98] = 1;cactus_sprite[4][22][99] = 1;cactus_sprite[4][23][13] = 1;cactus_sprite[4][23][14] = 1;cactus_sprite[4][23][15] = 1;cactus_sprite[4][23][16] = 1;cactus_sprite[4][23][17] = 1;cactus_sprite[4][23][18] = 1;cactus_sprite[4][23][19] = 1;cactus_sprite[4][23][20] = 1;cactus_sprite[4][23][21] = 1;cactus_sprite[4][23][22] = 1;cactus_sprite[4][23][23] = 1;cactus_sprite[4][23][24] = 1;cactus_sprite[4][23][25] = 1;cactus_sprite[4][23][26] = 1;cactus_sprite[4][23][27] = 1;cactus_sprite[4][23][28] = 1;cactus_sprite[4][23][29] = 1;cactus_sprite[4][23][30] = 1;cactus_sprite[4][23][31] = 1;cactus_sprite[4][23][32] = 1;cactus_sprite[4][23][33] = 1;cactus_sprite[4][23][34] = 1;cactus_sprite[4][23][35] = 1;cactus_sprite[4][23][36] = 1;cactus_sprite[4][23][37] = 1;cactus_sprite[4][23][38] = 1;cactus_sprite[4][23][39] = 1;cactus_sprite[4][23][40] = 1;cactus_sprite[4][23][41] = 1;cactus_sprite[4][23][42] = 1;cactus_sprite[4][23][43] = 1;cactus_sprite[4][23][44] = 1;cactus_sprite[4][23][45] = 1;cactus_sprite[4][23][46] = 1;cactus_sprite[4][23][47] = 1;cactus_sprite[4][23][48] = 1;cactus_sprite[4][23][49] = 1;cactus_sprite[4][23][50] = 1;cactus_sprite[4][23][51] = 1;cactus_sprite[4][23][52] = 1;cactus_sprite[4][23][53] = 1;cactus_sprite[4][23][54] = 1;cactus_sprite[4][23][55] = 1;cactus_sprite[4][23][56] = 1;cactus_sprite[4][23][57] = 1;cactus_sprite[4][23][58] = 1;cactus_sprite[4][23][59] = 1;cactus_sprite[4][23][60] = 1;cactus_sprite[4][23][61] = 1;cactus_sprite[4][23][62] = 1;cactus_sprite[4][23][63] = 1;cactus_sprite[4][23][64] = 1;cactus_sprite[4][23][65] = 1;cactus_sprite[4][23][66] = 1;cactus_sprite[4][23][67] = 1;cactus_sprite[4][23][68] = 1;cactus_sprite[4][23][69] = 1;cactus_sprite[4][23][70] = 1;cactus_sprite[4][23][71] = 1;cactus_sprite[4][23][72] = 1;cactus_sprite[4][23][73] = 1;cactus_sprite[4][23][74] = 1;cactus_sprite[4][23][75] = 1;cactus_sprite[4][23][76] = 1;cactus_sprite[4][23][77] = 1;cactus_sprite[4][23][78] = 1;cactus_sprite[4][23][79] = 1;cactus_sprite[4][23][80] = 1;cactus_sprite[4][23][81] = 1;cactus_sprite[4][23][82] = 1;cactus_sprite[4][23][83] = 1;cactus_sprite[4][23][84] = 1;cactus_sprite[4][23][85] = 1;cactus_sprite[4][23][86] = 1;cactus_sprite[4][23][87] = 1;cactus_sprite[4][23][88] = 1;cactus_sprite[4][23][89] = 1;cactus_sprite[4][23][90] = 1;cactus_sprite[4][23][91] = 1;cactus_sprite[4][23][92] = 1;cactus_sprite[4][23][93] = 1;cactus_sprite[4][23][94] = 1;cactus_sprite[4][23][95] = 1;cactus_sprite[4][23][96] = 1;cactus_sprite[4][23][97] = 1;cactus_sprite[4][23][98] = 1;cactus_sprite[4][23][99] = 1;cactus_sprite[4][24][41] = 1;cactus_sprite[4][24][42] = 1;cactus_sprite[4][24][43] = 1;cactus_sprite[4][24][44] = 1;cactus_sprite[4][24][45] = 1;cactus_sprite[4][24][46] = 1;cactus_sprite[4][25][41] = 1;cactus_sprite[4][25][42] = 1;cactus_sprite[4][25][43] = 1;cactus_sprite[4][25][44] = 1;cactus_sprite[4][25][45] = 1;cactus_sprite[4][25][46] = 1;cactus_sprite[4][26][41] = 1;cactus_sprite[4][26][42] = 1;cactus_sprite[4][26][43] = 1;cactus_sprite[4][26][44] = 1;cactus_sprite[4][26][45] = 1;cactus_sprite[4][26][46] = 1;cactus_sprite[4][27][41] = 1;cactus_sprite[4][27][42] = 1;cactus_sprite[4][27][43] = 1;cactus_sprite[4][27][44] = 1;cactus_sprite[4][27][45] = 1;cactus_sprite[4][27][46] = 1;cactus_sprite[4][28][41] = 1;cactus_sprite[4][28][42] = 1;cactus_sprite[4][28][43] = 1;cactus_sprite[4][28][44] = 1;cactus_sprite[4][28][45] = 1;cactus_sprite[4][28][46] = 1;cactus_sprite[4][29][41] = 1;cactus_sprite[4][29][42] = 1;cactus_sprite[4][29][43] = 1;cactus_sprite[4][29][44] = 1;cactus_sprite[4][29][45] = 1;cactus_sprite[4][29][46] = 1;cactus_sprite[4][30][23] = 1;cactus_sprite[4][30][24] = 1;cactus_sprite[4][30][25] = 1;cactus_sprite[4][30][26] = 1;cactus_sprite[4][30][27] = 1;cactus_sprite[4][30][28] = 1;cactus_sprite[4][30][29] = 1;cactus_sprite[4][30][30] = 1;cactus_sprite[4][30][31] = 1;cactus_sprite[4][30][32] = 1;cactus_sprite[4][30][33] = 1;cactus_sprite[4][30][34] = 1;cactus_sprite[4][30][35] = 1;cactus_sprite[4][30][36] = 1;cactus_sprite[4][30][37] = 1;cactus_sprite[4][30][38] = 1;cactus_sprite[4][30][39] = 1;cactus_sprite[4][30][40] = 1;cactus_sprite[4][30][41] = 1;cactus_sprite[4][30][42] = 1;cactus_sprite[4][30][43] = 1;cactus_sprite[4][30][44] = 1;cactus_sprite[4][30][45] = 1;cactus_sprite[4][30][46] = 1;cactus_sprite[4][31][23] = 1;cactus_sprite[4][31][24] = 1;cactus_sprite[4][31][25] = 1;cactus_sprite[4][31][26] = 1;cactus_sprite[4][31][27] = 1;cactus_sprite[4][31][28] = 1;cactus_sprite[4][31][29] = 1;cactus_sprite[4][31][30] = 1;cactus_sprite[4][31][31] = 1;cactus_sprite[4][31][32] = 1;cactus_sprite[4][31][33] = 1;cactus_sprite[4][31][34] = 1;cactus_sprite[4][31][35] = 1;cactus_sprite[4][31][36] = 1;cactus_sprite[4][31][37] = 1;cactus_sprite[4][31][38] = 1;cactus_sprite[4][31][39] = 1;cactus_sprite[4][31][40] = 1;cactus_sprite[4][31][41] = 1;cactus_sprite[4][31][42] = 1;cactus_sprite[4][31][43] = 1;cactus_sprite[4][31][44] = 1;cactus_sprite[4][31][45] = 1;cactus_sprite[4][31][46] = 1;cactus_sprite[4][32][21] = 1;cactus_sprite[4][32][22] = 1;cactus_sprite[4][32][23] = 1;cactus_sprite[4][32][24] = 1;cactus_sprite[4][32][25] = 1;cactus_sprite[4][32][26] = 1;cactus_sprite[4][32][27] = 1;cactus_sprite[4][32][28] = 1;cactus_sprite[4][32][29] = 1;cactus_sprite[4][32][30] = 1;cactus_sprite[4][32][31] = 1;cactus_sprite[4][32][32] = 1;cactus_sprite[4][32][33] = 1;cactus_sprite[4][32][34] = 1;cactus_sprite[4][32][35] = 1;cactus_sprite[4][32][36] = 1;cactus_sprite[4][32][37] = 1;cactus_sprite[4][32][38] = 1;cactus_sprite[4][32][39] = 1;cactus_sprite[4][32][40] = 1;cactus_sprite[4][32][41] = 1;cactus_sprite[4][32][42] = 1;cactus_sprite[4][32][43] = 1;cactus_sprite[4][32][44] = 1;cactus_sprite[4][33][21] = 1;cactus_sprite[4][33][22] = 1;cactus_sprite[4][33][23] = 1;cactus_sprite[4][33][24] = 1;cactus_sprite[4][33][25] = 1;cactus_sprite[4][33][26] = 1;cactus_sprite[4][33][27] = 1;cactus_sprite[4][33][28] = 1;cactus_sprite[4][33][29] = 1;cactus_sprite[4][33][30] = 1;cactus_sprite[4][33][31] = 1;cactus_sprite[4][33][32] = 1;cactus_sprite[4][33][33] = 1;cactus_sprite[4][33][34] = 1;cactus_sprite[4][33][35] = 1;cactus_sprite[4][33][36] = 1;cactus_sprite[4][33][37] = 1;cactus_sprite[4][33][38] = 1;cactus_sprite[4][33][39] = 1;cactus_sprite[4][33][40] = 1;cactus_sprite[4][33][41] = 1;cactus_sprite[4][33][42] = 1;cactus_sprite[4][33][43] = 1;cactus_sprite[4][33][44] = 1;cactus_sprite[4][34][23] = 1;cactus_sprite[4][34][24] = 1;cactus_sprite[4][34][25] = 1;cactus_sprite[4][34][26] = 1;cactus_sprite[4][34][27] = 1;cactus_sprite[4][34][28] = 1;cactus_sprite[4][34][29] = 1;cactus_sprite[4][34][30] = 1;cactus_sprite[4][34][31] = 1;cactus_sprite[4][34][32] = 1;cactus_sprite[4][34][33] = 1;cactus_sprite[4][34][34] = 1;cactus_sprite[4][34][35] = 1;cactus_sprite[4][34][36] = 1;cactus_sprite[4][34][37] = 1;cactus_sprite[4][34][38] = 1;cactus_sprite[4][34][39] = 1;cactus_sprite[4][34][40] = 1;cactus_sprite[4][34][41] = 1;cactus_sprite[4][34][42] = 1;cactus_sprite[4][35][23] = 1;cactus_sprite[4][35][24] = 1;cactus_sprite[4][35][25] = 1;cactus_sprite[4][35][26] = 1;cactus_sprite[4][35][27] = 1;cactus_sprite[4][35][28] = 1;cactus_sprite[4][35][29] = 1;cactus_sprite[4][35][30] = 1;cactus_sprite[4][35][31] = 1;cactus_sprite[4][35][32] = 1;cactus_sprite[4][35][33] = 1;cactus_sprite[4][35][34] = 1;cactus_sprite[4][35][35] = 1;cactus_sprite[4][35][36] = 1;cactus_sprite[4][35][37] = 1;cactus_sprite[4][35][38] = 1;cactus_sprite[4][35][39] = 1;cactus_sprite[4][35][40] = 1;cactus_sprite[4][35][41] = 1;cactus_sprite[4][35][42] = 1;
	cactus_sprite[5][2][20] = 1;cactus_sprite[5][2][21] = 1;cactus_sprite[5][2][22] = 1;cactus_sprite[5][2][23] = 1;cactus_sprite[5][2][24] = 1;cactus_sprite[5][2][25] = 1;cactus_sprite[5][2][26] = 1;cactus_sprite[5][2][27] = 1;cactus_sprite[5][2][28] = 1;cactus_sprite[5][2][29] = 1;cactus_sprite[5][2][30] = 1;cactus_sprite[5][2][31] = 1;cactus_sprite[5][2][32] = 1;cactus_sprite[5][2][33] = 1;cactus_sprite[5][2][34] = 1;cactus_sprite[5][2][35] = 1;cactus_sprite[5][2][36] = 1;cactus_sprite[5][2][37] = 1;cactus_sprite[5][2][38] = 1;cactus_sprite[5][2][39] = 1;cactus_sprite[5][2][40] = 1;cactus_sprite[5][2][41] = 1;cactus_sprite[5][2][42] = 1;cactus_sprite[5][2][43] = 1;cactus_sprite[5][2][44] = 1;cactus_sprite[5][2][45] = 1;cactus_sprite[5][2][46] = 1;cactus_sprite[5][2][47] = 1;cactus_sprite[5][2][48] = 1;cactus_sprite[5][2][49] = 1;cactus_sprite[5][3][20] = 1;cactus_sprite[5][3][21] = 1;cactus_sprite[5][3][22] = 1;cactus_sprite[5][3][23] = 1;cactus_sprite[5][3][24] = 1;cactus_sprite[5][3][25] = 1;cactus_sprite[5][3][26] = 1;cactus_sprite[5][3][27] = 1;cactus_sprite[5][3][28] = 1;cactus_sprite[5][3][29] = 1;cactus_sprite[5][3][30] = 1;cactus_sprite[5][3][31] = 1;cactus_sprite[5][3][32] = 1;cactus_sprite[5][3][33] = 1;cactus_sprite[5][3][34] = 1;cactus_sprite[5][3][35] = 1;cactus_sprite[5][3][36] = 1;cactus_sprite[5][3][37] = 1;cactus_sprite[5][3][38] = 1;cactus_sprite[5][3][39] = 1;cactus_sprite[5][3][40] = 1;cactus_sprite[5][3][41] = 1;cactus_sprite[5][3][42] = 1;cactus_sprite[5][3][43] = 1;cactus_sprite[5][3][44] = 1;cactus_sprite[5][3][45] = 1;cactus_sprite[5][3][46] = 1;cactus_sprite[5][3][47] = 1;cactus_sprite[5][3][48] = 1;cactus_sprite[5][3][49] = 1;cactus_sprite[5][4][18] = 1;cactus_sprite[5][4][19] = 1;cactus_sprite[5][4][20] = 1;cactus_sprite[5][4][21] = 1;cactus_sprite[5][4][22] = 1;cactus_sprite[5][4][23] = 1;cactus_sprite[5][4][24] = 1;cactus_sprite[5][4][25] = 1;cactus_sprite[5][4][26] = 1;cactus_sprite[5][4][27] = 1;cactus_sprite[5][4][28] = 1;cactus_sprite[5][4][29] = 1;cactus_sprite[5][4][30] = 1;cactus_sprite[5][4][31] = 1;cactus_sprite[5][4][32] = 1;cactus_sprite[5][4][33] = 1;cactus_sprite[5][4][34] = 1;cactus_sprite[5][4][35] = 1;cactus_sprite[5][4][36] = 1;cactus_sprite[5][4][37] = 1;cactus_sprite[5][4][38] = 1;cactus_sprite[5][4][39] = 1;cactus_sprite[5][4][40] = 1;cactus_sprite[5][4][41] = 1;cactus_sprite[5][4][42] = 1;cactus_sprite[5][4][43] = 1;cactus_sprite[5][4][44] = 1;cactus_sprite[5][4][45] = 1;cactus_sprite[5][4][46] = 1;cactus_sprite[5][4][47] = 1;cactus_sprite[5][4][48] = 1;cactus_sprite[5][4][49] = 1;cactus_sprite[5][4][50] = 1;cactus_sprite[5][4][51] = 1;cactus_sprite[5][5][18] = 1;cactus_sprite[5][5][19] = 1;cactus_sprite[5][5][20] = 1;cactus_sprite[5][5][21] = 1;cactus_sprite[5][5][22] = 1;cactus_sprite[5][5][23] = 1;cactus_sprite[5][5][24] = 1;cactus_sprite[5][5][25] = 1;cactus_sprite[5][5][26] = 1;cactus_sprite[5][5][27] = 1;cactus_sprite[5][5][28] = 1;cactus_sprite[5][5][29] = 1;cactus_sprite[5][5][30] = 1;cactus_sprite[5][5][31] = 1;cactus_sprite[5][5][32] = 1;cactus_sprite[5][5][33] = 1;cactus_sprite[5][5][34] = 1;cactus_sprite[5][5][35] = 1;cactus_sprite[5][5][36] = 1;cactus_sprite[5][5][37] = 1;cactus_sprite[5][5][38] = 1;cactus_sprite[5][5][39] = 1;cactus_sprite[5][5][40] = 1;cactus_sprite[5][5][41] = 1;cactus_sprite[5][5][42] = 1;cactus_sprite[5][5][43] = 1;cactus_sprite[5][5][44] = 1;cactus_sprite[5][5][45] = 1;cactus_sprite[5][5][46] = 1;cactus_sprite[5][5][47] = 1;cactus_sprite[5][5][48] = 1;cactus_sprite[5][5][49] = 1;cactus_sprite[5][5][50] = 1;cactus_sprite[5][5][51] = 1;cactus_sprite[5][6][18] = 1;cactus_sprite[5][6][19] = 1;cactus_sprite[5][6][20] = 1;cactus_sprite[5][6][21] = 1;cactus_sprite[5][6][22] = 1;cactus_sprite[5][6][23] = 1;cactus_sprite[5][6][24] = 1;cactus_sprite[5][6][25] = 1;cactus_sprite[5][6][26] = 1;cactus_sprite[5][6][27] = 1;cactus_sprite[5][6][28] = 1;cactus_sprite[5][6][29] = 1;cactus_sprite[5][6][30] = 1;cactus_sprite[5][6][31] = 1;cactus_sprite[5][6][32] = 1;cactus_sprite[5][6][33] = 1;cactus_sprite[5][6][34] = 1;cactus_sprite[5][6][35] = 1;cactus_sprite[5][6][36] = 1;cactus_sprite[5][6][37] = 1;cactus_sprite[5][6][38] = 1;cactus_sprite[5][6][39] = 1;cactus_sprite[5][6][40] = 1;cactus_sprite[5][6][41] = 1;cactus_sprite[5][6][42] = 1;cactus_sprite[5][6][43] = 1;cactus_sprite[5][6][44] = 1;cactus_sprite[5][6][45] = 1;cactus_sprite[5][6][46] = 1;cactus_sprite[5][6][47] = 1;cactus_sprite[5][6][48] = 1;cactus_sprite[5][6][49] = 1;cactus_sprite[5][6][50] = 1;cactus_sprite[5][6][51] = 1;cactus_sprite[5][6][52] = 1;cactus_sprite[5][6][53] = 1;cactus_sprite[5][7][18] = 1;cactus_sprite[5][7][19] = 1;cactus_sprite[5][7][20] = 1;cactus_sprite[5][7][21] = 1;cactus_sprite[5][7][22] = 1;cactus_sprite[5][7][23] = 1;cactus_sprite[5][7][24] = 1;cactus_sprite[5][7][25] = 1;cactus_sprite[5][7][26] = 1;cactus_sprite[5][7][27] = 1;cactus_sprite[5][7][28] = 1;cactus_sprite[5][7][29] = 1;cactus_sprite[5][7][30] = 1;cactus_sprite[5][7][31] = 1;cactus_sprite[5][7][32] = 1;cactus_sprite[5][7][33] = 1;cactus_sprite[5][7][34] = 1;cactus_sprite[5][7][35] = 1;cactus_sprite[5][7][36] = 1;cactus_sprite[5][7][37] = 1;cactus_sprite[5][7][38] = 1;cactus_sprite[5][7][39] = 1;cactus_sprite[5][7][40] = 1;cactus_sprite[5][7][41] = 1;cactus_sprite[5][7][42] = 1;cactus_sprite[5][7][43] = 1;cactus_sprite[5][7][44] = 1;cactus_sprite[5][7][45] = 1;cactus_sprite[5][7][46] = 1;cactus_sprite[5][7][47] = 1;cactus_sprite[5][7][48] = 1;cactus_sprite[5][7][49] = 1;cactus_sprite[5][7][50] = 1;cactus_sprite[5][7][51] = 1;cactus_sprite[5][7][52] = 1;cactus_sprite[5][7][53] = 1;cactus_sprite[5][8][18] = 1;cactus_sprite[5][8][19] = 1;cactus_sprite[5][8][20] = 1;cactus_sprite[5][8][21] = 1;cactus_sprite[5][8][22] = 1;cactus_sprite[5][8][23] = 1;cactus_sprite[5][8][24] = 1;cactus_sprite[5][8][25] = 1;cactus_sprite[5][8][26] = 1;cactus_sprite[5][8][27] = 1;cactus_sprite[5][8][28] = 1;cactus_sprite[5][8][29] = 1;cactus_sprite[5][8][30] = 1;cactus_sprite[5][8][31] = 1;cactus_sprite[5][8][32] = 1;cactus_sprite[5][8][33] = 1;cactus_sprite[5][8][34] = 1;cactus_sprite[5][8][35] = 1;cactus_sprite[5][8][36] = 1;cactus_sprite[5][8][37] = 1;cactus_sprite[5][8][38] = 1;cactus_sprite[5][8][39] = 1;cactus_sprite[5][8][40] = 1;cactus_sprite[5][8][41] = 1;cactus_sprite[5][8][42] = 1;cactus_sprite[5][8][43] = 1;cactus_sprite[5][8][44] = 1;cactus_sprite[5][8][45] = 1;cactus_sprite[5][8][46] = 1;cactus_sprite[5][8][47] = 1;cactus_sprite[5][8][48] = 1;cactus_sprite[5][8][49] = 1;cactus_sprite[5][8][50] = 1;cactus_sprite[5][8][51] = 1;cactus_sprite[5][8][52] = 1;cactus_sprite[5][8][53] = 1;cactus_sprite[5][8][54] = 1;cactus_sprite[5][8][55] = 1;cactus_sprite[5][9][18] = 1;cactus_sprite[5][9][19] = 1;cactus_sprite[5][9][20] = 1;cactus_sprite[5][9][21] = 1;cactus_sprite[5][9][22] = 1;cactus_sprite[5][9][23] = 1;cactus_sprite[5][9][24] = 1;cactus_sprite[5][9][25] = 1;cactus_sprite[5][9][26] = 1;cactus_sprite[5][9][27] = 1;cactus_sprite[5][9][28] = 1;cactus_sprite[5][9][29] = 1;cactus_sprite[5][9][30] = 1;cactus_sprite[5][9][31] = 1;cactus_sprite[5][9][32] = 1;cactus_sprite[5][9][33] = 1;cactus_sprite[5][9][34] = 1;cactus_sprite[5][9][35] = 1;cactus_sprite[5][9][36] = 1;cactus_sprite[5][9][37] = 1;cactus_sprite[5][9][38] = 1;cactus_sprite[5][9][39] = 1;cactus_sprite[5][9][40] = 1;cactus_sprite[5][9][41] = 1;cactus_sprite[5][9][42] = 1;cactus_sprite[5][9][43] = 1;cactus_sprite[5][9][44] = 1;cactus_sprite[5][9][45] = 1;cactus_sprite[5][9][46] = 1;cactus_sprite[5][9][47] = 1;cactus_sprite[5][9][48] = 1;cactus_sprite[5][9][49] = 1;cactus_sprite[5][9][50] = 1;cactus_sprite[5][9][51] = 1;cactus_sprite[5][9][52] = 1;cactus_sprite[5][9][53] = 1;cactus_sprite[5][9][54] = 1;cactus_sprite[5][9][55] = 1;cactus_sprite[5][10][20] = 1;cactus_sprite[5][10][21] = 1;cactus_sprite[5][10][22] = 1;cactus_sprite[5][10][23] = 1;cactus_sprite[5][10][24] = 1;cactus_sprite[5][10][25] = 1;cactus_sprite[5][10][26] = 1;cactus_sprite[5][10][27] = 1;cactus_sprite[5][10][28] = 1;cactus_sprite[5][10][29] = 1;cactus_sprite[5][10][30] = 1;cactus_sprite[5][10][31] = 1;cactus_sprite[5][10][32] = 1;cactus_sprite[5][10][33] = 1;cactus_sprite[5][10][34] = 1;cactus_sprite[5][10][35] = 1;cactus_sprite[5][10][36] = 1;cactus_sprite[5][10][37] = 1;cactus_sprite[5][10][38] = 1;cactus_sprite[5][10][39] = 1;cactus_sprite[5][10][40] = 1;cactus_sprite[5][10][41] = 1;cactus_sprite[5][10][42] = 1;cactus_sprite[5][10][43] = 1;cactus_sprite[5][10][44] = 1;cactus_sprite[5][10][45] = 1;cactus_sprite[5][10][46] = 1;cactus_sprite[5][10][47] = 1;cactus_sprite[5][10][48] = 1;cactus_sprite[5][10][49] = 1;cactus_sprite[5][10][50] = 1;cactus_sprite[5][10][51] = 1;cactus_sprite[5][10][52] = 1;cactus_sprite[5][10][53] = 1;cactus_sprite[5][10][54] = 1;cactus_sprite[5][10][55] = 1;cactus_sprite[5][11][20] = 1;cactus_sprite[5][11][21] = 1;cactus_sprite[5][11][22] = 1;cactus_sprite[5][11][23] = 1;cactus_sprite[5][11][24] = 1;cactus_sprite[5][11][25] = 1;cactus_sprite[5][11][26] = 1;cactus_sprite[5][11][27] = 1;cactus_sprite[5][11][28] = 1;cactus_sprite[5][11][29] = 1;cactus_sprite[5][11][30] = 1;cactus_sprite[5][11][31] = 1;cactus_sprite[5][11][32] = 1;cactus_sprite[5][11][33] = 1;cactus_sprite[5][11][34] = 1;cactus_sprite[5][11][35] = 1;cactus_sprite[5][11][36] = 1;cactus_sprite[5][11][37] = 1;cactus_sprite[5][11][38] = 1;cactus_sprite[5][11][39] = 1;cactus_sprite[5][11][40] = 1;cactus_sprite[5][11][41] = 1;cactus_sprite[5][11][42] = 1;cactus_sprite[5][11][43] = 1;cactus_sprite[5][11][44] = 1;cactus_sprite[5][11][45] = 1;cactus_sprite[5][11][46] = 1;cactus_sprite[5][11][47] = 1;cactus_sprite[5][11][48] = 1;cactus_sprite[5][11][49] = 1;cactus_sprite[5][11][50] = 1;cactus_sprite[5][11][51] = 1;cactus_sprite[5][11][52] = 1;cactus_sprite[5][11][53] = 1;cactus_sprite[5][11][54] = 1;cactus_sprite[5][11][55] = 1;cactus_sprite[5][12][46] = 1;cactus_sprite[5][12][47] = 1;cactus_sprite[5][12][48] = 1;cactus_sprite[5][12][49] = 1;cactus_sprite[5][12][50] = 1;cactus_sprite[5][12][51] = 1;cactus_sprite[5][12][52] = 1;cactus_sprite[5][12][53] = 1;cactus_sprite[5][12][54] = 1;cactus_sprite[5][12][55] = 1;cactus_sprite[5][13][46] = 1;cactus_sprite[5][13][47] = 1;cactus_sprite[5][13][48] = 1;cactus_sprite[5][13][49] = 1;cactus_sprite[5][13][50] = 1;cactus_sprite[5][13][51] = 1;cactus_sprite[5][13][52] = 1;cactus_sprite[5][13][53] = 1;cactus_sprite[5][13][54] = 1;cactus_sprite[5][13][55] = 1;cactus_sprite[5][14][46] = 1;cactus_sprite[5][14][47] = 1;cactus_sprite[5][14][48] = 1;cactus_sprite[5][14][49] = 1;cactus_sprite[5][14][50] = 1;cactus_sprite[5][14][51] = 1;cactus_sprite[5][14][52] = 1;cactus_sprite[5][14][53] = 1;cactus_sprite[5][14][54] = 1;cactus_sprite[5][14][55] = 1;cactus_sprite[5][14][98] = 1;cactus_sprite[5][14][99] = 1;cactus_sprite[5][15][46] = 1;cactus_sprite[5][15][47] = 1;cactus_sprite[5][15][48] = 1;cactus_sprite[5][15][49] = 1;cactus_sprite[5][15][50] = 1;cactus_sprite[5][15][51] = 1;cactus_sprite[5][15][52] = 1;cactus_sprite[5][15][53] = 1;cactus_sprite[5][15][54] = 1;cactus_sprite[5][15][55] = 1;cactus_sprite[5][15][98] = 1;cactus_sprite[5][15][99] = 1;cactus_sprite[5][16][46] = 1;cactus_sprite[5][16][47] = 1;cactus_sprite[5][16][48] = 1;cactus_sprite[5][16][49] = 1;cactus_sprite[5][16][50] = 1;cactus_sprite[5][16][51] = 1;cactus_sprite[5][16][52] = 1;cactus_sprite[5][16][53] = 1;cactus_sprite[5][16][54] = 1;cactus_sprite[5][16][55] = 1;cactus_sprite[5][16][98] = 1;cactus_sprite[5][16][99] = 1;cactus_sprite[5][17][46] = 1;cactus_sprite[5][17][47] = 1;cactus_sprite[5][17][48] = 1;cactus_sprite[5][17][49] = 1;cactus_sprite[5][17][50] = 1;cactus_sprite[5][17][51] = 1;cactus_sprite[5][17][52] = 1;cactus_sprite[5][17][53] = 1;cactus_sprite[5][17][54] = 1;cactus_sprite[5][17][55] = 1;cactus_sprite[5][17][98] = 1;cactus_sprite[5][17][99] = 1;cactus_sprite[5][18][8] = 1;cactus_sprite[5][18][9] = 1;cactus_sprite[5][18][10] = 1;cactus_sprite[5][18][11] = 1;cactus_sprite[5][18][12] = 1;cactus_sprite[5][18][13] = 1;cactus_sprite[5][18][14] = 1;cactus_sprite[5][18][15] = 1;cactus_sprite[5][18][16] = 1;cactus_sprite[5][18][17] = 1;cactus_sprite[5][18][18] = 1;cactus_sprite[5][18][19] = 1;cactus_sprite[5][18][20] = 1;cactus_sprite[5][18][21] = 1;cactus_sprite[5][18][22] = 1;cactus_sprite[5][18][23] = 1;cactus_sprite[5][18][24] = 1;cactus_sprite[5][18][25] = 1;cactus_sprite[5][18][26] = 1;cactus_sprite[5][18][27] = 1;cactus_sprite[5][18][28] = 1;cactus_sprite[5][18][29] = 1;cactus_sprite[5][18][30] = 1;cactus_sprite[5][18][31] = 1;cactus_sprite[5][18][32] = 1;cactus_sprite[5][18][33] = 1;cactus_sprite[5][18][34] = 1;cactus_sprite[5][18][35] = 1;cactus_sprite[5][18][36] = 1;cactus_sprite[5][18][37] = 1;cactus_sprite[5][18][38] = 1;cactus_sprite[5][18][39] = 1;cactus_sprite[5][18][40] = 1;cactus_sprite[5][18][41] = 1;cactus_sprite[5][18][42] = 1;cactus_sprite[5][18][43] = 1;cactus_sprite[5][18][44] = 1;cactus_sprite[5][18][45] = 1;cactus_sprite[5][18][46] = 1;cactus_sprite[5][18][47] = 1;cactus_sprite[5][18][48] = 1;cactus_sprite[5][18][49] = 1;cactus_sprite[5][18][50] = 1;cactus_sprite[5][18][51] = 1;cactus_sprite[5][18][52] = 1;cactus_sprite[5][18][53] = 1;cactus_sprite[5][18][54] = 1;cactus_sprite[5][18][55] = 1;cactus_sprite[5][18][56] = 1;cactus_sprite[5][18][57] = 1;cactus_sprite[5][18][58] = 1;cactus_sprite[5][18][59] = 1;cactus_sprite[5][18][60] = 1;cactus_sprite[5][18][61] = 1;cactus_sprite[5][18][62] = 1;cactus_sprite[5][18][63] = 1;cactus_sprite[5][18][64] = 1;cactus_sprite[5][18][65] = 1;cactus_sprite[5][18][66] = 1;cactus_sprite[5][18][67] = 1;cactus_sprite[5][18][68] = 1;cactus_sprite[5][18][69] = 1;cactus_sprite[5][18][70] = 1;cactus_sprite[5][18][71] = 1;cactus_sprite[5][18][72] = 1;cactus_sprite[5][18][73] = 1;cactus_sprite[5][18][74] = 1;cactus_sprite[5][18][75] = 1;cactus_sprite[5][18][76] = 1;cactus_sprite[5][18][77] = 1;cactus_sprite[5][18][78] = 1;cactus_sprite[5][18][79] = 1;cactus_sprite[5][18][80] = 1;cactus_sprite[5][18][81] = 1;cactus_sprite[5][18][82] = 1;cactus_sprite[5][18][83] = 1;cactus_sprite[5][18][84] = 1;cactus_sprite[5][18][85] = 1;cactus_sprite[5][18][86] = 1;cactus_sprite[5][18][87] = 1;cactus_sprite[5][18][88] = 1;cactus_sprite[5][18][89] = 1;cactus_sprite[5][18][90] = 1;cactus_sprite[5][18][91] = 1;cactus_sprite[5][18][92] = 1;cactus_sprite[5][18][93] = 1;cactus_sprite[5][18][94] = 1;cactus_sprite[5][18][95] = 1;cactus_sprite[5][18][96] = 1;cactus_sprite[5][18][97] = 1;cactus_sprite[5][18][98] = 1;cactus_sprite[5][18][99] = 1;cactus_sprite[5][19][8] = 1;cactus_sprite[5][19][9] = 1;cactus_sprite[5][19][10] = 1;cactus_sprite[5][19][11] = 1;cactus_sprite[5][19][12] = 1;cactus_sprite[5][19][13] = 1;cactus_sprite[5][19][14] = 1;cactus_sprite[5][19][15] = 1;cactus_sprite[5][19][16] = 1;cactus_sprite[5][19][17] = 1;cactus_sprite[5][19][18] = 1;cactus_sprite[5][19][19] = 1;cactus_sprite[5][19][20] = 1;cactus_sprite[5][19][21] = 1;cactus_sprite[5][19][22] = 1;cactus_sprite[5][19][23] = 1;cactus_sprite[5][19][24] = 1;cactus_sprite[5][19][25] = 1;cactus_sprite[5][19][26] = 1;cactus_sprite[5][19][27] = 1;cactus_sprite[5][19][28] = 1;cactus_sprite[5][19][29] = 1;cactus_sprite[5][19][30] = 1;cactus_sprite[5][19][31] = 1;cactus_sprite[5][19][32] = 1;cactus_sprite[5][19][33] = 1;cactus_sprite[5][19][34] = 1;cactus_sprite[5][19][35] = 1;cactus_sprite[5][19][36] = 1;cactus_sprite[5][19][37] = 1;cactus_sprite[5][19][38] = 1;cactus_sprite[5][19][39] = 1;cactus_sprite[5][19][40] = 1;cactus_sprite[5][19][41] = 1;cactus_sprite[5][19][42] = 1;cactus_sprite[5][19][43] = 1;cactus_sprite[5][19][44] = 1;cactus_sprite[5][19][45] = 1;cactus_sprite[5][19][46] = 1;cactus_sprite[5][19][47] = 1;cactus_sprite[5][19][48] = 1;cactus_sprite[5][19][49] = 1;cactus_sprite[5][19][50] = 1;cactus_sprite[5][19][51] = 1;cactus_sprite[5][19][52] = 1;cactus_sprite[5][19][53] = 1;cactus_sprite[5][19][54] = 1;cactus_sprite[5][19][55] = 1;cactus_sprite[5][19][56] = 1;cactus_sprite[5][19][57] = 1;cactus_sprite[5][19][58] = 1;cactus_sprite[5][19][59] = 1;cactus_sprite[5][19][60] = 1;cactus_sprite[5][19][61] = 1;cactus_sprite[5][19][62] = 1;cactus_sprite[5][19][63] = 1;cactus_sprite[5][19][64] = 1;cactus_sprite[5][19][65] = 1;cactus_sprite[5][19][66] = 1;cactus_sprite[5][19][67] = 1;cactus_sprite[5][19][68] = 1;cactus_sprite[5][19][69] = 1;cactus_sprite[5][19][70] = 1;cactus_sprite[5][19][71] = 1;cactus_sprite[5][19][72] = 1;cactus_sprite[5][19][73] = 1;cactus_sprite[5][19][74] = 1;cactus_sprite[5][19][75] = 1;cactus_sprite[5][19][76] = 1;cactus_sprite[5][19][77] = 1;cactus_sprite[5][19][78] = 1;cactus_sprite[5][19][79] = 1;cactus_sprite[5][19][80] = 1;cactus_sprite[5][19][81] = 1;cactus_sprite[5][19][82] = 1;cactus_sprite[5][19][83] = 1;cactus_sprite[5][19][84] = 1;cactus_sprite[5][19][85] = 1;cactus_sprite[5][19][86] = 1;cactus_sprite[5][19][87] = 1;cactus_sprite[5][19][88] = 1;cactus_sprite[5][19][89] = 1;cactus_sprite[5][19][90] = 1;cactus_sprite[5][19][91] = 1;cactus_sprite[5][19][92] = 1;cactus_sprite[5][19][93] = 1;cactus_sprite[5][19][94] = 1;cactus_sprite[5][19][95] = 1;cactus_sprite[5][19][96] = 1;cactus_sprite[5][19][97] = 1;cactus_sprite[5][19][98] = 1;cactus_sprite[5][19][99] = 1;cactus_sprite[5][20][6] = 1;cactus_sprite[5][20][7] = 1;cactus_sprite[5][20][8] = 1;cactus_sprite[5][20][9] = 1;cactus_sprite[5][20][10] = 1;cactus_sprite[5][20][11] = 1;cactus_sprite[5][20][12] = 1;cactus_sprite[5][20][13] = 1;cactus_sprite[5][20][14] = 1;cactus_sprite[5][20][15] = 1;cactus_sprite[5][20][16] = 1;cactus_sprite[5][20][17] = 1;cactus_sprite[5][20][18] = 1;cactus_sprite[5][20][19] = 1;cactus_sprite[5][20][20] = 1;cactus_sprite[5][20][21] = 1;cactus_sprite[5][20][22] = 1;cactus_sprite[5][20][23] = 1;cactus_sprite[5][20][24] = 1;cactus_sprite[5][20][25] = 1;cactus_sprite[5][20][26] = 1;cactus_sprite[5][20][27] = 1;cactus_sprite[5][20][28] = 1;cactus_sprite[5][20][29] = 1;cactus_sprite[5][20][30] = 1;cactus_sprite[5][20][31] = 1;cactus_sprite[5][20][32] = 1;cactus_sprite[5][20][33] = 1;cactus_sprite[5][20][34] = 1;cactus_sprite[5][20][35] = 1;cactus_sprite[5][20][36] = 1;cactus_sprite[5][20][37] = 1;cactus_sprite[5][20][38] = 1;cactus_sprite[5][20][39] = 1;cactus_sprite[5][20][40] = 1;cactus_sprite[5][20][41] = 1;cactus_sprite[5][20][42] = 1;cactus_sprite[5][20][43] = 1;cactus_sprite[5][20][44] = 1;cactus_sprite[5][20][45] = 1;cactus_sprite[5][20][46] = 1;cactus_sprite[5][20][47] = 1;cactus_sprite[5][20][48] = 1;cactus_sprite[5][20][49] = 1;cactus_sprite[5][20][50] = 1;cactus_sprite[5][20][51] = 1;cactus_sprite[5][20][52] = 1;cactus_sprite[5][20][53] = 1;cactus_sprite[5][20][54] = 1;cactus_sprite[5][20][55] = 1;cactus_sprite[5][20][56] = 1;cactus_sprite[5][20][57] = 1;cactus_sprite[5][20][58] = 1;cactus_sprite[5][20][59] = 1;cactus_sprite[5][20][60] = 1;cactus_sprite[5][20][61] = 1;cactus_sprite[5][20][62] = 1;cactus_sprite[5][20][63] = 1;cactus_sprite[5][20][64] = 1;cactus_sprite[5][20][65] = 1;cactus_sprite[5][20][66] = 1;cactus_sprite[5][20][67] = 1;cactus_sprite[5][20][68] = 1;cactus_sprite[5][20][69] = 1;cactus_sprite[5][20][70] = 1;cactus_sprite[5][20][71] = 1;cactus_sprite[5][20][72] = 1;cactus_sprite[5][20][73] = 1;cactus_sprite[5][20][74] = 1;cactus_sprite[5][20][75] = 1;cactus_sprite[5][20][76] = 1;cactus_sprite[5][20][77] = 1;cactus_sprite[5][20][78] = 1;cactus_sprite[5][20][79] = 1;cactus_sprite[5][20][80] = 1;cactus_sprite[5][20][81] = 1;cactus_sprite[5][20][82] = 1;cactus_sprite[5][20][83] = 1;cactus_sprite[5][20][84] = 1;cactus_sprite[5][20][85] = 1;cactus_sprite[5][20][86] = 1;cactus_sprite[5][20][87] = 1;cactus_sprite[5][20][88] = 1;cactus_sprite[5][20][89] = 1;cactus_sprite[5][20][90] = 1;cactus_sprite[5][20][91] = 1;cactus_sprite[5][20][92] = 1;cactus_sprite[5][20][93] = 1;cactus_sprite[5][20][94] = 1;cactus_sprite[5][20][95] = 1;cactus_sprite[5][20][96] = 1;cactus_sprite[5][20][97] = 1;cactus_sprite[5][20][98] = 1;cactus_sprite[5][20][99] = 1;cactus_sprite[5][21][6] = 1;cactus_sprite[5][21][7] = 1;cactus_sprite[5][21][8] = 1;cactus_sprite[5][21][9] = 1;cactus_sprite[5][21][10] = 1;cactus_sprite[5][21][11] = 1;cactus_sprite[5][21][12] = 1;cactus_sprite[5][21][13] = 1;cactus_sprite[5][21][14] = 1;cactus_sprite[5][21][15] = 1;cactus_sprite[5][21][16] = 1;cactus_sprite[5][21][17] = 1;cactus_sprite[5][21][18] = 1;cactus_sprite[5][21][19] = 1;cactus_sprite[5][21][20] = 1;cactus_sprite[5][21][21] = 1;cactus_sprite[5][21][22] = 1;cactus_sprite[5][21][23] = 1;cactus_sprite[5][21][24] = 1;cactus_sprite[5][21][25] = 1;cactus_sprite[5][21][26] = 1;cactus_sprite[5][21][27] = 1;cactus_sprite[5][21][28] = 1;cactus_sprite[5][21][29] = 1;cactus_sprite[5][21][30] = 1;cactus_sprite[5][21][31] = 1;cactus_sprite[5][21][32] = 1;cactus_sprite[5][21][33] = 1;cactus_sprite[5][21][34] = 1;cactus_sprite[5][21][35] = 1;cactus_sprite[5][21][36] = 1;cactus_sprite[5][21][37] = 1;cactus_sprite[5][21][38] = 1;cactus_sprite[5][21][39] = 1;cactus_sprite[5][21][40] = 1;cactus_sprite[5][21][41] = 1;cactus_sprite[5][21][42] = 1;cactus_sprite[5][21][43] = 1;cactus_sprite[5][21][44] = 1;cactus_sprite[5][21][45] = 1;cactus_sprite[5][21][46] = 1;cactus_sprite[5][21][47] = 1;cactus_sprite[5][21][48] = 1;cactus_sprite[5][21][49] = 1;cactus_sprite[5][21][50] = 1;cactus_sprite[5][21][51] = 1;cactus_sprite[5][21][52] = 1;cactus_sprite[5][21][53] = 1;cactus_sprite[5][21][54] = 1;cactus_sprite[5][21][55] = 1;cactus_sprite[5][21][56] = 1;cactus_sprite[5][21][57] = 1;cactus_sprite[5][21][58] = 1;cactus_sprite[5][21][59] = 1;cactus_sprite[5][21][60] = 1;cactus_sprite[5][21][61] = 1;cactus_sprite[5][21][62] = 1;cactus_sprite[5][21][63] = 1;cactus_sprite[5][21][64] = 1;cactus_sprite[5][21][65] = 1;cactus_sprite[5][21][66] = 1;cactus_sprite[5][21][67] = 1;cactus_sprite[5][21][68] = 1;cactus_sprite[5][21][69] = 1;cactus_sprite[5][21][70] = 1;cactus_sprite[5][21][71] = 1;cactus_sprite[5][21][72] = 1;cactus_sprite[5][21][73] = 1;cactus_sprite[5][21][74] = 1;cactus_sprite[5][21][75] = 1;cactus_sprite[5][21][76] = 1;cactus_sprite[5][21][77] = 1;cactus_sprite[5][21][78] = 1;cactus_sprite[5][21][79] = 1;cactus_sprite[5][21][80] = 1;cactus_sprite[5][21][81] = 1;cactus_sprite[5][21][82] = 1;cactus_sprite[5][21][83] = 1;cactus_sprite[5][21][84] = 1;cactus_sprite[5][21][85] = 1;cactus_sprite[5][21][86] = 1;cactus_sprite[5][21][87] = 1;cactus_sprite[5][21][88] = 1;cactus_sprite[5][21][89] = 1;cactus_sprite[5][21][90] = 1;cactus_sprite[5][21][91] = 1;cactus_sprite[5][21][92] = 1;cactus_sprite[5][21][93] = 1;cactus_sprite[5][21][94] = 1;cactus_sprite[5][21][95] = 1;cactus_sprite[5][21][96] = 1;cactus_sprite[5][21][97] = 1;cactus_sprite[5][21][98] = 1;cactus_sprite[5][21][99] = 1;cactus_sprite[5][22][6] = 1;cactus_sprite[5][22][7] = 1;cactus_sprite[5][22][8] = 1;cactus_sprite[5][22][9] = 1;cactus_sprite[5][22][10] = 1;cactus_sprite[5][22][11] = 1;cactus_sprite[5][22][12] = 1;cactus_sprite[5][22][13] = 1;cactus_sprite[5][22][14] = 1;cactus_sprite[5][22][15] = 1;cactus_sprite[5][22][16] = 1;cactus_sprite[5][22][17] = 1;cactus_sprite[5][22][18] = 1;cactus_sprite[5][22][19] = 1;cactus_sprite[5][22][20] = 1;cactus_sprite[5][22][21] = 1;cactus_sprite[5][22][22] = 1;cactus_sprite[5][22][23] = 1;cactus_sprite[5][22][24] = 1;cactus_sprite[5][22][25] = 1;cactus_sprite[5][22][26] = 1;cactus_sprite[5][22][27] = 1;cactus_sprite[5][22][28] = 1;cactus_sprite[5][22][29] = 1;cactus_sprite[5][22][30] = 1;cactus_sprite[5][22][31] = 1;cactus_sprite[5][22][32] = 1;cactus_sprite[5][22][33] = 1;cactus_sprite[5][22][34] = 1;cactus_sprite[5][22][35] = 1;cactus_sprite[5][22][36] = 1;cactus_sprite[5][22][37] = 1;cactus_sprite[5][22][38] = 1;cactus_sprite[5][22][39] = 1;cactus_sprite[5][22][40] = 1;cactus_sprite[5][22][41] = 1;cactus_sprite[5][22][42] = 1;cactus_sprite[5][22][43] = 1;cactus_sprite[5][22][44] = 1;cactus_sprite[5][22][45] = 1;cactus_sprite[5][22][46] = 1;cactus_sprite[5][22][47] = 1;cactus_sprite[5][22][48] = 1;cactus_sprite[5][22][49] = 1;cactus_sprite[5][22][50] = 1;cactus_sprite[5][22][51] = 1;cactus_sprite[5][22][52] = 1;cactus_sprite[5][22][53] = 1;cactus_sprite[5][22][54] = 1;cactus_sprite[5][22][55] = 1;cactus_sprite[5][22][56] = 1;cactus_sprite[5][22][57] = 1;cactus_sprite[5][22][58] = 1;cactus_sprite[5][22][59] = 1;cactus_sprite[5][22][60] = 1;cactus_sprite[5][22][61] = 1;cactus_sprite[5][22][62] = 1;cactus_sprite[5][22][63] = 1;cactus_sprite[5][22][64] = 1;cactus_sprite[5][22][65] = 1;cactus_sprite[5][22][66] = 1;cactus_sprite[5][22][67] = 1;cactus_sprite[5][22][68] = 1;cactus_sprite[5][22][69] = 1;cactus_sprite[5][22][70] = 1;cactus_sprite[5][22][71] = 1;cactus_sprite[5][22][72] = 1;cactus_sprite[5][22][73] = 1;cactus_sprite[5][22][74] = 1;cactus_sprite[5][22][75] = 1;cactus_sprite[5][22][76] = 1;cactus_sprite[5][22][77] = 1;cactus_sprite[5][22][78] = 1;cactus_sprite[5][22][79] = 1;cactus_sprite[5][22][80] = 1;cactus_sprite[5][22][81] = 1;cactus_sprite[5][22][82] = 1;cactus_sprite[5][22][83] = 1;cactus_sprite[5][22][84] = 1;cactus_sprite[5][22][85] = 1;cactus_sprite[5][22][86] = 1;cactus_sprite[5][22][87] = 1;cactus_sprite[5][22][88] = 1;cactus_sprite[5][22][89] = 1;cactus_sprite[5][22][90] = 1;cactus_sprite[5][22][91] = 1;cactus_sprite[5][22][92] = 1;cactus_sprite[5][22][93] = 1;cactus_sprite[5][22][94] = 1;cactus_sprite[5][22][95] = 1;cactus_sprite[5][22][96] = 1;cactus_sprite[5][22][97] = 1;cactus_sprite[5][22][98] = 1;cactus_sprite[5][22][99] = 1;cactus_sprite[5][23][6] = 1;cactus_sprite[5][23][7] = 1;cactus_sprite[5][23][8] = 1;cactus_sprite[5][23][9] = 1;cactus_sprite[5][23][10] = 1;cactus_sprite[5][23][11] = 1;cactus_sprite[5][23][12] = 1;cactus_sprite[5][23][13] = 1;cactus_sprite[5][23][14] = 1;cactus_sprite[5][23][15] = 1;cactus_sprite[5][23][16] = 1;cactus_sprite[5][23][17] = 1;cactus_sprite[5][23][18] = 1;cactus_sprite[5][23][19] = 1;cactus_sprite[5][23][20] = 1;cactus_sprite[5][23][21] = 1;cactus_sprite[5][23][22] = 1;cactus_sprite[5][23][23] = 1;cactus_sprite[5][23][24] = 1;cactus_sprite[5][23][25] = 1;cactus_sprite[5][23][26] = 1;cactus_sprite[5][23][27] = 1;cactus_sprite[5][23][28] = 1;cactus_sprite[5][23][29] = 1;cactus_sprite[5][23][30] = 1;cactus_sprite[5][23][31] = 1;cactus_sprite[5][23][32] = 1;cactus_sprite[5][23][33] = 1;cactus_sprite[5][23][34] = 1;cactus_sprite[5][23][35] = 1;cactus_sprite[5][23][36] = 1;cactus_sprite[5][23][37] = 1;cactus_sprite[5][23][38] = 1;cactus_sprite[5][23][39] = 1;cactus_sprite[5][23][40] = 1;cactus_sprite[5][23][41] = 1;cactus_sprite[5][23][42] = 1;cactus_sprite[5][23][43] = 1;cactus_sprite[5][23][44] = 1;cactus_sprite[5][23][45] = 1;cactus_sprite[5][23][46] = 1;cactus_sprite[5][23][47] = 1;cactus_sprite[5][23][48] = 1;cactus_sprite[5][23][49] = 1;cactus_sprite[5][23][50] = 1;cactus_sprite[5][23][51] = 1;cactus_sprite[5][23][52] = 1;cactus_sprite[5][23][53] = 1;cactus_sprite[5][23][54] = 1;cactus_sprite[5][23][55] = 1;cactus_sprite[5][23][56] = 1;cactus_sprite[5][23][57] = 1;cactus_sprite[5][23][58] = 1;cactus_sprite[5][23][59] = 1;cactus_sprite[5][23][60] = 1;cactus_sprite[5][23][61] = 1;cactus_sprite[5][23][62] = 1;cactus_sprite[5][23][63] = 1;cactus_sprite[5][23][64] = 1;cactus_sprite[5][23][65] = 1;cactus_sprite[5][23][66] = 1;cactus_sprite[5][23][67] = 1;cactus_sprite[5][23][68] = 1;cactus_sprite[5][23][69] = 1;cactus_sprite[5][23][70] = 1;cactus_sprite[5][23][71] = 1;cactus_sprite[5][23][72] = 1;cactus_sprite[5][23][73] = 1;cactus_sprite[5][23][74] = 1;cactus_sprite[5][23][75] = 1;cactus_sprite[5][23][76] = 1;cactus_sprite[5][23][77] = 1;cactus_sprite[5][23][78] = 1;cactus_sprite[5][23][79] = 1;cactus_sprite[5][23][80] = 1;cactus_sprite[5][23][81] = 1;cactus_sprite[5][23][82] = 1;cactus_sprite[5][23][83] = 1;cactus_sprite[5][23][84] = 1;cactus_sprite[5][23][85] = 1;cactus_sprite[5][23][86] = 1;cactus_sprite[5][23][87] = 1;cactus_sprite[5][23][88] = 1;cactus_sprite[5][23][89] = 1;cactus_sprite[5][23][90] = 1;cactus_sprite[5][23][91] = 1;cactus_sprite[5][23][92] = 1;cactus_sprite[5][23][93] = 1;cactus_sprite[5][23][94] = 1;cactus_sprite[5][23][95] = 1;cactus_sprite[5][23][96] = 1;cactus_sprite[5][23][97] = 1;cactus_sprite[5][23][98] = 1;cactus_sprite[5][23][99] = 1;cactus_sprite[5][24][6] = 1;cactus_sprite[5][24][7] = 1;cactus_sprite[5][24][8] = 1;cactus_sprite[5][24][9] = 1;cactus_sprite[5][24][10] = 1;cactus_sprite[5][24][11] = 1;cactus_sprite[5][24][12] = 1;cactus_sprite[5][24][13] = 1;cactus_sprite[5][24][14] = 1;cactus_sprite[5][24][15] = 1;cactus_sprite[5][24][16] = 1;cactus_sprite[5][24][17] = 1;cactus_sprite[5][24][18] = 1;cactus_sprite[5][24][19] = 1;cactus_sprite[5][24][20] = 1;cactus_sprite[5][24][21] = 1;cactus_sprite[5][24][22] = 1;cactus_sprite[5][24][23] = 1;cactus_sprite[5][24][24] = 1;cactus_sprite[5][24][25] = 1;cactus_sprite[5][24][26] = 1;cactus_sprite[5][24][27] = 1;cactus_sprite[5][24][28] = 1;cactus_sprite[5][24][29] = 1;cactus_sprite[5][24][30] = 1;cactus_sprite[5][24][31] = 1;cactus_sprite[5][24][32] = 1;cactus_sprite[5][24][33] = 1;cactus_sprite[5][24][34] = 1;cactus_sprite[5][24][35] = 1;cactus_sprite[5][24][36] = 1;cactus_sprite[5][24][37] = 1;cactus_sprite[5][24][38] = 1;cactus_sprite[5][24][39] = 1;cactus_sprite[5][24][40] = 1;cactus_sprite[5][24][41] = 1;cactus_sprite[5][24][42] = 1;cactus_sprite[5][24][43] = 1;cactus_sprite[5][24][44] = 1;cactus_sprite[5][24][45] = 1;cactus_sprite[5][24][46] = 1;cactus_sprite[5][24][47] = 1;cactus_sprite[5][24][48] = 1;cactus_sprite[5][24][49] = 1;cactus_sprite[5][24][50] = 1;cactus_sprite[5][24][51] = 1;cactus_sprite[5][24][52] = 1;cactus_sprite[5][24][53] = 1;cactus_sprite[5][24][54] = 1;cactus_sprite[5][24][55] = 1;cactus_sprite[5][24][56] = 1;cactus_sprite[5][24][57] = 1;cactus_sprite[5][24][58] = 1;cactus_sprite[5][24][59] = 1;cactus_sprite[5][24][60] = 1;cactus_sprite[5][24][61] = 1;cactus_sprite[5][24][62] = 1;cactus_sprite[5][24][63] = 1;cactus_sprite[5][24][64] = 1;cactus_sprite[5][24][65] = 1;cactus_sprite[5][24][66] = 1;cactus_sprite[5][24][67] = 1;cactus_sprite[5][24][68] = 1;cactus_sprite[5][24][69] = 1;cactus_sprite[5][24][70] = 1;cactus_sprite[5][24][71] = 1;cactus_sprite[5][24][72] = 1;cactus_sprite[5][24][73] = 1;cactus_sprite[5][24][74] = 1;cactus_sprite[5][24][75] = 1;cactus_sprite[5][24][76] = 1;cactus_sprite[5][24][77] = 1;cactus_sprite[5][24][78] = 1;cactus_sprite[5][24][79] = 1;cactus_sprite[5][24][80] = 1;cactus_sprite[5][24][81] = 1;cactus_sprite[5][24][82] = 1;cactus_sprite[5][24][83] = 1;cactus_sprite[5][24][84] = 1;cactus_sprite[5][24][85] = 1;cactus_sprite[5][24][86] = 1;cactus_sprite[5][24][87] = 1;cactus_sprite[5][24][88] = 1;cactus_sprite[5][24][89] = 1;cactus_sprite[5][24][90] = 1;cactus_sprite[5][24][91] = 1;cactus_sprite[5][24][92] = 1;cactus_sprite[5][24][93] = 1;cactus_sprite[5][24][94] = 1;cactus_sprite[5][24][95] = 1;cactus_sprite[5][24][96] = 1;cactus_sprite[5][24][97] = 1;cactus_sprite[5][24][98] = 1;cactus_sprite[5][24][99] = 1;cactus_sprite[5][25][6] = 1;cactus_sprite[5][25][7] = 1;cactus_sprite[5][25][8] = 1;cactus_sprite[5][25][9] = 1;cactus_sprite[5][25][10] = 1;cactus_sprite[5][25][11] = 1;cactus_sprite[5][25][12] = 1;cactus_sprite[5][25][13] = 1;cactus_sprite[5][25][14] = 1;cactus_sprite[5][25][15] = 1;cactus_sprite[5][25][16] = 1;cactus_sprite[5][25][17] = 1;cactus_sprite[5][25][18] = 1;cactus_sprite[5][25][19] = 1;cactus_sprite[5][25][20] = 1;cactus_sprite[5][25][21] = 1;cactus_sprite[5][25][22] = 1;cactus_sprite[5][25][23] = 1;cactus_sprite[5][25][24] = 1;cactus_sprite[5][25][25] = 1;cactus_sprite[5][25][26] = 1;cactus_sprite[5][25][27] = 1;cactus_sprite[5][25][28] = 1;cactus_sprite[5][25][29] = 1;cactus_sprite[5][25][30] = 1;cactus_sprite[5][25][31] = 1;cactus_sprite[5][25][32] = 1;cactus_sprite[5][25][33] = 1;cactus_sprite[5][25][34] = 1;cactus_sprite[5][25][35] = 1;cactus_sprite[5][25][36] = 1;cactus_sprite[5][25][37] = 1;cactus_sprite[5][25][38] = 1;cactus_sprite[5][25][39] = 1;cactus_sprite[5][25][40] = 1;cactus_sprite[5][25][41] = 1;cactus_sprite[5][25][42] = 1;cactus_sprite[5][25][43] = 1;cactus_sprite[5][25][44] = 1;cactus_sprite[5][25][45] = 1;cactus_sprite[5][25][46] = 1;cactus_sprite[5][25][47] = 1;cactus_sprite[5][25][48] = 1;cactus_sprite[5][25][49] = 1;cactus_sprite[5][25][50] = 1;cactus_sprite[5][25][51] = 1;cactus_sprite[5][25][52] = 1;cactus_sprite[5][25][53] = 1;cactus_sprite[5][25][54] = 1;cactus_sprite[5][25][55] = 1;cactus_sprite[5][25][56] = 1;cactus_sprite[5][25][57] = 1;cactus_sprite[5][25][58] = 1;cactus_sprite[5][25][59] = 1;cactus_sprite[5][25][60] = 1;cactus_sprite[5][25][61] = 1;cactus_sprite[5][25][62] = 1;cactus_sprite[5][25][63] = 1;cactus_sprite[5][25][64] = 1;cactus_sprite[5][25][65] = 1;cactus_sprite[5][25][66] = 1;cactus_sprite[5][25][67] = 1;cactus_sprite[5][25][68] = 1;cactus_sprite[5][25][69] = 1;cactus_sprite[5][25][70] = 1;cactus_sprite[5][25][71] = 1;cactus_sprite[5][25][72] = 1;cactus_sprite[5][25][73] = 1;cactus_sprite[5][25][74] = 1;cactus_sprite[5][25][75] = 1;cactus_sprite[5][25][76] = 1;cactus_sprite[5][25][77] = 1;cactus_sprite[5][25][78] = 1;cactus_sprite[5][25][79] = 1;cactus_sprite[5][25][80] = 1;cactus_sprite[5][25][81] = 1;cactus_sprite[5][25][82] = 1;cactus_sprite[5][25][83] = 1;cactus_sprite[5][25][84] = 1;cactus_sprite[5][25][85] = 1;cactus_sprite[5][25][86] = 1;cactus_sprite[5][25][87] = 1;cactus_sprite[5][25][88] = 1;cactus_sprite[5][25][89] = 1;cactus_sprite[5][25][90] = 1;cactus_sprite[5][25][91] = 1;cactus_sprite[5][25][92] = 1;cactus_sprite[5][25][93] = 1;cactus_sprite[5][25][94] = 1;cactus_sprite[5][25][95] = 1;cactus_sprite[5][25][96] = 1;cactus_sprite[5][25][97] = 1;cactus_sprite[5][25][98] = 1;cactus_sprite[5][25][99] = 1;cactus_sprite[5][26][6] = 1;cactus_sprite[5][26][7] = 1;cactus_sprite[5][26][8] = 1;cactus_sprite[5][26][9] = 1;cactus_sprite[5][26][10] = 1;cactus_sprite[5][26][11] = 1;cactus_sprite[5][26][12] = 1;cactus_sprite[5][26][13] = 1;cactus_sprite[5][26][14] = 1;cactus_sprite[5][26][15] = 1;cactus_sprite[5][26][16] = 1;cactus_sprite[5][26][17] = 1;cactus_sprite[5][26][18] = 1;cactus_sprite[5][26][19] = 1;cactus_sprite[5][26][20] = 1;cactus_sprite[5][26][21] = 1;cactus_sprite[5][26][22] = 1;cactus_sprite[5][26][23] = 1;cactus_sprite[5][26][24] = 1;cactus_sprite[5][26][25] = 1;cactus_sprite[5][26][26] = 1;cactus_sprite[5][26][27] = 1;cactus_sprite[5][26][28] = 1;cactus_sprite[5][26][29] = 1;cactus_sprite[5][26][30] = 1;cactus_sprite[5][26][31] = 1;cactus_sprite[5][26][32] = 1;cactus_sprite[5][26][33] = 1;cactus_sprite[5][26][34] = 1;cactus_sprite[5][26][35] = 1;cactus_sprite[5][26][36] = 1;cactus_sprite[5][26][37] = 1;cactus_sprite[5][26][38] = 1;cactus_sprite[5][26][39] = 1;cactus_sprite[5][26][40] = 1;cactus_sprite[5][26][41] = 1;cactus_sprite[5][26][42] = 1;cactus_sprite[5][26][43] = 1;cactus_sprite[5][26][44] = 1;cactus_sprite[5][26][45] = 1;cactus_sprite[5][26][46] = 1;cactus_sprite[5][26][47] = 1;cactus_sprite[5][26][48] = 1;cactus_sprite[5][26][49] = 1;cactus_sprite[5][26][50] = 1;cactus_sprite[5][26][51] = 1;cactus_sprite[5][26][52] = 1;cactus_sprite[5][26][53] = 1;cactus_sprite[5][26][54] = 1;cactus_sprite[5][26][55] = 1;cactus_sprite[5][26][56] = 1;cactus_sprite[5][26][57] = 1;cactus_sprite[5][26][58] = 1;cactus_sprite[5][26][59] = 1;cactus_sprite[5][26][60] = 1;cactus_sprite[5][26][61] = 1;cactus_sprite[5][26][62] = 1;cactus_sprite[5][26][63] = 1;cactus_sprite[5][26][64] = 1;cactus_sprite[5][26][65] = 1;cactus_sprite[5][26][66] = 1;cactus_sprite[5][26][67] = 1;cactus_sprite[5][26][68] = 1;cactus_sprite[5][26][69] = 1;cactus_sprite[5][26][70] = 1;cactus_sprite[5][26][71] = 1;cactus_sprite[5][26][72] = 1;cactus_sprite[5][26][73] = 1;cactus_sprite[5][26][74] = 1;cactus_sprite[5][26][75] = 1;cactus_sprite[5][26][76] = 1;cactus_sprite[5][26][77] = 1;cactus_sprite[5][26][78] = 1;cactus_sprite[5][26][79] = 1;cactus_sprite[5][26][80] = 1;cactus_sprite[5][26][81] = 1;cactus_sprite[5][26][82] = 1;cactus_sprite[5][26][83] = 1;cactus_sprite[5][26][84] = 1;cactus_sprite[5][26][85] = 1;cactus_sprite[5][26][86] = 1;cactus_sprite[5][26][87] = 1;cactus_sprite[5][26][88] = 1;cactus_sprite[5][26][89] = 1;cactus_sprite[5][26][90] = 1;cactus_sprite[5][26][91] = 1;cactus_sprite[5][26][92] = 1;cactus_sprite[5][26][93] = 1;cactus_sprite[5][26][94] = 1;cactus_sprite[5][26][95] = 1;cactus_sprite[5][26][96] = 1;cactus_sprite[5][26][97] = 1;cactus_sprite[5][26][98] = 1;cactus_sprite[5][26][99] = 1;cactus_sprite[5][27][6] = 1;cactus_sprite[5][27][7] = 1;cactus_sprite[5][27][8] = 1;cactus_sprite[5][27][9] = 1;cactus_sprite[5][27][10] = 1;cactus_sprite[5][27][11] = 1;cactus_sprite[5][27][12] = 1;cactus_sprite[5][27][13] = 1;cactus_sprite[5][27][14] = 1;cactus_sprite[5][27][15] = 1;cactus_sprite[5][27][16] = 1;cactus_sprite[5][27][17] = 1;cactus_sprite[5][27][18] = 1;cactus_sprite[5][27][19] = 1;cactus_sprite[5][27][20] = 1;cactus_sprite[5][27][21] = 1;cactus_sprite[5][27][22] = 1;cactus_sprite[5][27][23] = 1;cactus_sprite[5][27][24] = 1;cactus_sprite[5][27][25] = 1;cactus_sprite[5][27][26] = 1;cactus_sprite[5][27][27] = 1;cactus_sprite[5][27][28] = 1;cactus_sprite[5][27][29] = 1;cactus_sprite[5][27][30] = 1;cactus_sprite[5][27][31] = 1;cactus_sprite[5][27][32] = 1;cactus_sprite[5][27][33] = 1;cactus_sprite[5][27][34] = 1;cactus_sprite[5][27][35] = 1;cactus_sprite[5][27][36] = 1;cactus_sprite[5][27][37] = 1;cactus_sprite[5][27][38] = 1;cactus_sprite[5][27][39] = 1;cactus_sprite[5][27][40] = 1;cactus_sprite[5][27][41] = 1;cactus_sprite[5][27][42] = 1;cactus_sprite[5][27][43] = 1;cactus_sprite[5][27][44] = 1;cactus_sprite[5][27][45] = 1;cactus_sprite[5][27][46] = 1;cactus_sprite[5][27][47] = 1;cactus_sprite[5][27][48] = 1;cactus_sprite[5][27][49] = 1;cactus_sprite[5][27][50] = 1;cactus_sprite[5][27][51] = 1;cactus_sprite[5][27][52] = 1;cactus_sprite[5][27][53] = 1;cactus_sprite[5][27][54] = 1;cactus_sprite[5][27][55] = 1;cactus_sprite[5][27][56] = 1;cactus_sprite[5][27][57] = 1;cactus_sprite[5][27][58] = 1;cactus_sprite[5][27][59] = 1;cactus_sprite[5][27][60] = 1;cactus_sprite[5][27][61] = 1;cactus_sprite[5][27][62] = 1;cactus_sprite[5][27][63] = 1;cactus_sprite[5][27][64] = 1;cactus_sprite[5][27][65] = 1;cactus_sprite[5][27][66] = 1;cactus_sprite[5][27][67] = 1;cactus_sprite[5][27][68] = 1;cactus_sprite[5][27][69] = 1;cactus_sprite[5][27][70] = 1;cactus_sprite[5][27][71] = 1;cactus_sprite[5][27][72] = 1;cactus_sprite[5][27][73] = 1;cactus_sprite[5][27][74] = 1;cactus_sprite[5][27][75] = 1;cactus_sprite[5][27][76] = 1;cactus_sprite[5][27][77] = 1;cactus_sprite[5][27][78] = 1;cactus_sprite[5][27][79] = 1;cactus_sprite[5][27][80] = 1;cactus_sprite[5][27][81] = 1;cactus_sprite[5][27][82] = 1;cactus_sprite[5][27][83] = 1;cactus_sprite[5][27][84] = 1;cactus_sprite[5][27][85] = 1;cactus_sprite[5][27][86] = 1;cactus_sprite[5][27][87] = 1;cactus_sprite[5][27][88] = 1;cactus_sprite[5][27][89] = 1;cactus_sprite[5][27][90] = 1;cactus_sprite[5][27][91] = 1;cactus_sprite[5][27][92] = 1;cactus_sprite[5][27][93] = 1;cactus_sprite[5][27][94] = 1;cactus_sprite[5][27][95] = 1;cactus_sprite[5][27][96] = 1;cactus_sprite[5][27][97] = 1;cactus_sprite[5][27][98] = 1;cactus_sprite[5][27][99] = 1;cactus_sprite[5][28][6] = 1;cactus_sprite[5][28][7] = 1;cactus_sprite[5][28][8] = 1;cactus_sprite[5][28][9] = 1;cactus_sprite[5][28][10] = 1;cactus_sprite[5][28][11] = 1;cactus_sprite[5][28][12] = 1;cactus_sprite[5][28][13] = 1;cactus_sprite[5][28][14] = 1;cactus_sprite[5][28][15] = 1;cactus_sprite[5][28][16] = 1;cactus_sprite[5][28][17] = 1;cactus_sprite[5][28][18] = 1;cactus_sprite[5][28][19] = 1;cactus_sprite[5][28][20] = 1;cactus_sprite[5][28][21] = 1;cactus_sprite[5][28][22] = 1;cactus_sprite[5][28][23] = 1;cactus_sprite[5][28][24] = 1;cactus_sprite[5][28][25] = 1;cactus_sprite[5][28][26] = 1;cactus_sprite[5][28][27] = 1;cactus_sprite[5][28][28] = 1;cactus_sprite[5][28][29] = 1;cactus_sprite[5][28][30] = 1;cactus_sprite[5][28][31] = 1;cactus_sprite[5][28][32] = 1;cactus_sprite[5][28][33] = 1;cactus_sprite[5][28][34] = 1;cactus_sprite[5][28][35] = 1;cactus_sprite[5][28][36] = 1;cactus_sprite[5][28][37] = 1;cactus_sprite[5][28][38] = 1;cactus_sprite[5][28][39] = 1;cactus_sprite[5][28][40] = 1;cactus_sprite[5][28][41] = 1;cactus_sprite[5][28][42] = 1;cactus_sprite[5][28][43] = 1;cactus_sprite[5][28][44] = 1;cactus_sprite[5][28][45] = 1;cactus_sprite[5][28][46] = 1;cactus_sprite[5][28][47] = 1;cactus_sprite[5][28][48] = 1;cactus_sprite[5][28][49] = 1;cactus_sprite[5][28][50] = 1;cactus_sprite[5][28][51] = 1;cactus_sprite[5][28][52] = 1;cactus_sprite[5][28][53] = 1;cactus_sprite[5][28][54] = 1;cactus_sprite[5][28][55] = 1;cactus_sprite[5][28][56] = 1;cactus_sprite[5][28][57] = 1;cactus_sprite[5][28][58] = 1;cactus_sprite[5][28][59] = 1;cactus_sprite[5][28][60] = 1;cactus_sprite[5][28][61] = 1;cactus_sprite[5][28][62] = 1;cactus_sprite[5][28][63] = 1;cactus_sprite[5][28][64] = 1;cactus_sprite[5][28][65] = 1;cactus_sprite[5][28][66] = 1;cactus_sprite[5][28][67] = 1;cactus_sprite[5][28][68] = 1;cactus_sprite[5][28][69] = 1;cactus_sprite[5][28][70] = 1;cactus_sprite[5][28][71] = 1;cactus_sprite[5][28][72] = 1;cactus_sprite[5][28][73] = 1;cactus_sprite[5][28][74] = 1;cactus_sprite[5][28][75] = 1;cactus_sprite[5][28][76] = 1;cactus_sprite[5][28][77] = 1;cactus_sprite[5][28][78] = 1;cactus_sprite[5][28][79] = 1;cactus_sprite[5][28][80] = 1;cactus_sprite[5][28][81] = 1;cactus_sprite[5][28][82] = 1;cactus_sprite[5][28][83] = 1;cactus_sprite[5][28][84] = 1;cactus_sprite[5][28][85] = 1;cactus_sprite[5][28][86] = 1;cactus_sprite[5][28][87] = 1;cactus_sprite[5][28][88] = 1;cactus_sprite[5][28][89] = 1;cactus_sprite[5][28][90] = 1;cactus_sprite[5][28][91] = 1;cactus_sprite[5][28][92] = 1;cactus_sprite[5][28][93] = 1;cactus_sprite[5][28][94] = 1;cactus_sprite[5][28][95] = 1;cactus_sprite[5][28][96] = 1;cactus_sprite[5][28][97] = 1;cactus_sprite[5][28][98] = 1;cactus_sprite[5][28][99] = 1;cactus_sprite[5][29][6] = 1;cactus_sprite[5][29][7] = 1;cactus_sprite[5][29][8] = 1;cactus_sprite[5][29][9] = 1;cactus_sprite[5][29][10] = 1;cactus_sprite[5][29][11] = 1;cactus_sprite[5][29][12] = 1;cactus_sprite[5][29][13] = 1;cactus_sprite[5][29][14] = 1;cactus_sprite[5][29][15] = 1;cactus_sprite[5][29][16] = 1;cactus_sprite[5][29][17] = 1;cactus_sprite[5][29][18] = 1;cactus_sprite[5][29][19] = 1;cactus_sprite[5][29][20] = 1;cactus_sprite[5][29][21] = 1;cactus_sprite[5][29][22] = 1;cactus_sprite[5][29][23] = 1;cactus_sprite[5][29][24] = 1;cactus_sprite[5][29][25] = 1;cactus_sprite[5][29][26] = 1;cactus_sprite[5][29][27] = 1;cactus_sprite[5][29][28] = 1;cactus_sprite[5][29][29] = 1;cactus_sprite[5][29][30] = 1;cactus_sprite[5][29][31] = 1;cactus_sprite[5][29][32] = 1;cactus_sprite[5][29][33] = 1;cactus_sprite[5][29][34] = 1;cactus_sprite[5][29][35] = 1;cactus_sprite[5][29][36] = 1;cactus_sprite[5][29][37] = 1;cactus_sprite[5][29][38] = 1;cactus_sprite[5][29][39] = 1;cactus_sprite[5][29][40] = 1;cactus_sprite[5][29][41] = 1;cactus_sprite[5][29][42] = 1;cactus_sprite[5][29][43] = 1;cactus_sprite[5][29][44] = 1;cactus_sprite[5][29][45] = 1;cactus_sprite[5][29][46] = 1;cactus_sprite[5][29][47] = 1;cactus_sprite[5][29][48] = 1;cactus_sprite[5][29][49] = 1;cactus_sprite[5][29][50] = 1;cactus_sprite[5][29][51] = 1;cactus_sprite[5][29][52] = 1;cactus_sprite[5][29][53] = 1;cactus_sprite[5][29][54] = 1;cactus_sprite[5][29][55] = 1;cactus_sprite[5][29][56] = 1;cactus_sprite[5][29][57] = 1;cactus_sprite[5][29][58] = 1;cactus_sprite[5][29][59] = 1;cactus_sprite[5][29][60] = 1;cactus_sprite[5][29][61] = 1;cactus_sprite[5][29][62] = 1;cactus_sprite[5][29][63] = 1;cactus_sprite[5][29][64] = 1;cactus_sprite[5][29][65] = 1;cactus_sprite[5][29][66] = 1;cactus_sprite[5][29][67] = 1;cactus_sprite[5][29][68] = 1;cactus_sprite[5][29][69] = 1;cactus_sprite[5][29][70] = 1;cactus_sprite[5][29][71] = 1;cactus_sprite[5][29][72] = 1;cactus_sprite[5][29][73] = 1;cactus_sprite[5][29][74] = 1;cactus_sprite[5][29][75] = 1;cactus_sprite[5][29][76] = 1;cactus_sprite[5][29][77] = 1;cactus_sprite[5][29][78] = 1;cactus_sprite[5][29][79] = 1;cactus_sprite[5][29][80] = 1;cactus_sprite[5][29][81] = 1;cactus_sprite[5][29][82] = 1;cactus_sprite[5][29][83] = 1;cactus_sprite[5][29][84] = 1;cactus_sprite[5][29][85] = 1;cactus_sprite[5][29][86] = 1;cactus_sprite[5][29][87] = 1;cactus_sprite[5][29][88] = 1;cactus_sprite[5][29][89] = 1;cactus_sprite[5][29][90] = 1;cactus_sprite[5][29][91] = 1;cactus_sprite[5][29][92] = 1;cactus_sprite[5][29][93] = 1;cactus_sprite[5][29][94] = 1;cactus_sprite[5][29][95] = 1;cactus_sprite[5][29][96] = 1;cactus_sprite[5][29][97] = 1;cactus_sprite[5][29][98] = 1;cactus_sprite[5][29][99] = 1;cactus_sprite[5][30][8] = 1;cactus_sprite[5][30][9] = 1;cactus_sprite[5][30][10] = 1;cactus_sprite[5][30][11] = 1;cactus_sprite[5][30][12] = 1;cactus_sprite[5][30][13] = 1;cactus_sprite[5][30][14] = 1;cactus_sprite[5][30][15] = 1;cactus_sprite[5][30][16] = 1;cactus_sprite[5][30][17] = 1;cactus_sprite[5][30][18] = 1;cactus_sprite[5][30][19] = 1;cactus_sprite[5][30][20] = 1;cactus_sprite[5][30][21] = 1;cactus_sprite[5][30][22] = 1;cactus_sprite[5][30][23] = 1;cactus_sprite[5][30][24] = 1;cactus_sprite[5][30][25] = 1;cactus_sprite[5][30][26] = 1;cactus_sprite[5][30][27] = 1;cactus_sprite[5][30][28] = 1;cactus_sprite[5][30][29] = 1;cactus_sprite[5][30][30] = 1;cactus_sprite[5][30][31] = 1;cactus_sprite[5][30][32] = 1;cactus_sprite[5][30][33] = 1;cactus_sprite[5][30][34] = 1;cactus_sprite[5][30][35] = 1;cactus_sprite[5][30][36] = 1;cactus_sprite[5][30][37] = 1;cactus_sprite[5][30][38] = 1;cactus_sprite[5][30][39] = 1;cactus_sprite[5][30][40] = 1;cactus_sprite[5][30][41] = 1;cactus_sprite[5][30][42] = 1;cactus_sprite[5][30][43] = 1;cactus_sprite[5][30][44] = 1;cactus_sprite[5][30][45] = 1;cactus_sprite[5][30][46] = 1;cactus_sprite[5][30][47] = 1;cactus_sprite[5][30][48] = 1;cactus_sprite[5][30][49] = 1;cactus_sprite[5][30][50] = 1;cactus_sprite[5][30][51] = 1;cactus_sprite[5][30][52] = 1;cactus_sprite[5][30][53] = 1;cactus_sprite[5][30][54] = 1;cactus_sprite[5][30][55] = 1;cactus_sprite[5][30][56] = 1;cactus_sprite[5][30][57] = 1;cactus_sprite[5][30][58] = 1;cactus_sprite[5][30][59] = 1;cactus_sprite[5][30][60] = 1;cactus_sprite[5][30][61] = 1;cactus_sprite[5][30][62] = 1;cactus_sprite[5][30][63] = 1;cactus_sprite[5][30][64] = 1;cactus_sprite[5][30][65] = 1;cactus_sprite[5][30][66] = 1;cactus_sprite[5][30][67] = 1;cactus_sprite[5][30][68] = 1;cactus_sprite[5][30][69] = 1;cactus_sprite[5][30][70] = 1;cactus_sprite[5][30][71] = 1;cactus_sprite[5][30][72] = 1;cactus_sprite[5][30][73] = 1;cactus_sprite[5][30][74] = 1;cactus_sprite[5][30][75] = 1;cactus_sprite[5][30][76] = 1;cactus_sprite[5][30][77] = 1;cactus_sprite[5][30][78] = 1;cactus_sprite[5][30][79] = 1;cactus_sprite[5][30][80] = 1;cactus_sprite[5][30][81] = 1;cactus_sprite[5][30][82] = 1;cactus_sprite[5][30][83] = 1;cactus_sprite[5][30][84] = 1;cactus_sprite[5][30][85] = 1;cactus_sprite[5][30][86] = 1;cactus_sprite[5][30][87] = 1;cactus_sprite[5][30][88] = 1;cactus_sprite[5][30][89] = 1;cactus_sprite[5][30][90] = 1;cactus_sprite[5][30][91] = 1;cactus_sprite[5][30][92] = 1;cactus_sprite[5][30][93] = 1;cactus_sprite[5][30][94] = 1;cactus_sprite[5][30][95] = 1;cactus_sprite[5][30][96] = 1;cactus_sprite[5][30][97] = 1;cactus_sprite[5][30][98] = 1;cactus_sprite[5][30][99] = 1;cactus_sprite[5][31][8] = 1;cactus_sprite[5][31][9] = 1;cactus_sprite[5][31][10] = 1;cactus_sprite[5][31][11] = 1;cactus_sprite[5][31][12] = 1;cactus_sprite[5][31][13] = 1;cactus_sprite[5][31][14] = 1;cactus_sprite[5][31][15] = 1;cactus_sprite[5][31][16] = 1;cactus_sprite[5][31][17] = 1;cactus_sprite[5][31][18] = 1;cactus_sprite[5][31][19] = 1;cactus_sprite[5][31][20] = 1;cactus_sprite[5][31][21] = 1;cactus_sprite[5][31][22] = 1;cactus_sprite[5][31][23] = 1;cactus_sprite[5][31][24] = 1;cactus_sprite[5][31][25] = 1;cactus_sprite[5][31][26] = 1;cactus_sprite[5][31][27] = 1;cactus_sprite[5][31][28] = 1;cactus_sprite[5][31][29] = 1;cactus_sprite[5][31][30] = 1;cactus_sprite[5][31][31] = 1;cactus_sprite[5][31][32] = 1;cactus_sprite[5][31][33] = 1;cactus_sprite[5][31][34] = 1;cactus_sprite[5][31][35] = 1;cactus_sprite[5][31][36] = 1;cactus_sprite[5][31][37] = 1;cactus_sprite[5][31][38] = 1;cactus_sprite[5][31][39] = 1;cactus_sprite[5][31][40] = 1;cactus_sprite[5][31][41] = 1;cactus_sprite[5][31][42] = 1;cactus_sprite[5][31][43] = 1;cactus_sprite[5][31][44] = 1;cactus_sprite[5][31][45] = 1;cactus_sprite[5][31][46] = 1;cactus_sprite[5][31][47] = 1;cactus_sprite[5][31][48] = 1;cactus_sprite[5][31][49] = 1;cactus_sprite[5][31][50] = 1;cactus_sprite[5][31][51] = 1;cactus_sprite[5][31][52] = 1;cactus_sprite[5][31][53] = 1;cactus_sprite[5][31][54] = 1;cactus_sprite[5][31][55] = 1;cactus_sprite[5][31][56] = 1;cactus_sprite[5][31][57] = 1;cactus_sprite[5][31][58] = 1;cactus_sprite[5][31][59] = 1;cactus_sprite[5][31][60] = 1;cactus_sprite[5][31][61] = 1;cactus_sprite[5][31][62] = 1;cactus_sprite[5][31][63] = 1;cactus_sprite[5][31][64] = 1;cactus_sprite[5][31][65] = 1;cactus_sprite[5][31][66] = 1;cactus_sprite[5][31][67] = 1;cactus_sprite[5][31][68] = 1;cactus_sprite[5][31][69] = 1;cactus_sprite[5][31][70] = 1;cactus_sprite[5][31][71] = 1;cactus_sprite[5][31][72] = 1;cactus_sprite[5][31][73] = 1;cactus_sprite[5][31][74] = 1;cactus_sprite[5][31][75] = 1;cactus_sprite[5][31][76] = 1;cactus_sprite[5][31][77] = 1;cactus_sprite[5][31][78] = 1;cactus_sprite[5][31][79] = 1;cactus_sprite[5][31][80] = 1;cactus_sprite[5][31][81] = 1;cactus_sprite[5][31][82] = 1;cactus_sprite[5][31][83] = 1;cactus_sprite[5][31][84] = 1;cactus_sprite[5][31][85] = 1;cactus_sprite[5][31][86] = 1;cactus_sprite[5][31][87] = 1;cactus_sprite[5][31][88] = 1;cactus_sprite[5][31][89] = 1;cactus_sprite[5][31][90] = 1;cactus_sprite[5][31][91] = 1;cactus_sprite[5][31][92] = 1;cactus_sprite[5][31][93] = 1;cactus_sprite[5][31][94] = 1;cactus_sprite[5][31][95] = 1;cactus_sprite[5][31][96] = 1;cactus_sprite[5][31][97] = 1;cactus_sprite[5][31][98] = 1;cactus_sprite[5][31][99] = 1;cactus_sprite[5][32][60] = 1;cactus_sprite[5][32][61] = 1;cactus_sprite[5][32][62] = 1;cactus_sprite[5][32][63] = 1;cactus_sprite[5][32][64] = 1;cactus_sprite[5][32][65] = 1;cactus_sprite[5][33][60] = 1;cactus_sprite[5][33][61] = 1;cactus_sprite[5][33][62] = 1;cactus_sprite[5][33][63] = 1;cactus_sprite[5][33][64] = 1;cactus_sprite[5][33][65] = 1;cactus_sprite[5][34][60] = 1;cactus_sprite[5][34][61] = 1;cactus_sprite[5][34][62] = 1;cactus_sprite[5][34][63] = 1;cactus_sprite[5][34][64] = 1;cactus_sprite[5][34][65] = 1;cactus_sprite[5][35][60] = 1;cactus_sprite[5][35][61] = 1;cactus_sprite[5][35][62] = 1;cactus_sprite[5][35][63] = 1;cactus_sprite[5][35][64] = 1;cactus_sprite[5][35][65] = 1;cactus_sprite[5][36][60] = 1;cactus_sprite[5][36][61] = 1;cactus_sprite[5][36][62] = 1;cactus_sprite[5][36][63] = 1;cactus_sprite[5][36][64] = 1;cactus_sprite[5][36][65] = 1;cactus_sprite[5][36][97] = 1;cactus_sprite[5][37][60] = 1;cactus_sprite[5][37][61] = 1;cactus_sprite[5][37][62] = 1;cactus_sprite[5][37][63] = 1;cactus_sprite[5][37][64] = 1;cactus_sprite[5][37][65] = 1;cactus_sprite[5][38][30] = 1;cactus_sprite[5][38][31] = 1;cactus_sprite[5][38][32] = 1;cactus_sprite[5][38][33] = 1;cactus_sprite[5][38][34] = 1;cactus_sprite[5][38][35] = 1;cactus_sprite[5][38][36] = 1;cactus_sprite[5][38][37] = 1;cactus_sprite[5][38][38] = 1;cactus_sprite[5][38][39] = 1;cactus_sprite[5][38][40] = 1;cactus_sprite[5][38][41] = 1;cactus_sprite[5][38][42] = 1;cactus_sprite[5][38][43] = 1;cactus_sprite[5][38][44] = 1;cactus_sprite[5][38][45] = 1;cactus_sprite[5][38][46] = 1;cactus_sprite[5][38][47] = 1;cactus_sprite[5][38][48] = 1;cactus_sprite[5][38][49] = 1;cactus_sprite[5][38][50] = 1;cactus_sprite[5][38][51] = 1;cactus_sprite[5][38][52] = 1;cactus_sprite[5][38][53] = 1;cactus_sprite[5][38][54] = 1;cactus_sprite[5][38][55] = 1;cactus_sprite[5][38][56] = 1;cactus_sprite[5][38][57] = 1;cactus_sprite[5][38][58] = 1;cactus_sprite[5][38][59] = 1;cactus_sprite[5][38][60] = 1;cactus_sprite[5][38][61] = 1;cactus_sprite[5][38][62] = 1;cactus_sprite[5][38][63] = 1;cactus_sprite[5][38][64] = 1;cactus_sprite[5][38][65] = 1;cactus_sprite[5][39][30] = 1;cactus_sprite[5][39][31] = 1;cactus_sprite[5][39][32] = 1;cactus_sprite[5][39][33] = 1;cactus_sprite[5][39][34] = 1;cactus_sprite[5][39][35] = 1;cactus_sprite[5][39][36] = 1;cactus_sprite[5][39][37] = 1;cactus_sprite[5][39][38] = 1;cactus_sprite[5][39][39] = 1;cactus_sprite[5][39][40] = 1;cactus_sprite[5][39][41] = 1;cactus_sprite[5][39][42] = 1;cactus_sprite[5][39][43] = 1;cactus_sprite[5][39][44] = 1;cactus_sprite[5][39][45] = 1;cactus_sprite[5][39][46] = 1;cactus_sprite[5][39][47] = 1;cactus_sprite[5][39][48] = 1;cactus_sprite[5][39][49] = 1;cactus_sprite[5][39][50] = 1;cactus_sprite[5][39][51] = 1;cactus_sprite[5][39][52] = 1;cactus_sprite[5][39][53] = 1;cactus_sprite[5][39][54] = 1;cactus_sprite[5][39][55] = 1;cactus_sprite[5][39][56] = 1;cactus_sprite[5][39][57] = 1;cactus_sprite[5][39][58] = 1;cactus_sprite[5][39][59] = 1;cactus_sprite[5][39][60] = 1;cactus_sprite[5][39][61] = 1;cactus_sprite[5][39][62] = 1;cactus_sprite[5][39][63] = 1;cactus_sprite[5][39][64] = 1;cactus_sprite[5][39][65] = 1;cactus_sprite[5][40][28] = 1;cactus_sprite[5][40][29] = 1;cactus_sprite[5][40][30] = 1;cactus_sprite[5][40][31] = 1;cactus_sprite[5][40][32] = 1;cactus_sprite[5][40][33] = 1;cactus_sprite[5][40][34] = 1;cactus_sprite[5][40][35] = 1;cactus_sprite[5][40][36] = 1;cactus_sprite[5][40][37] = 1;cactus_sprite[5][40][38] = 1;cactus_sprite[5][40][39] = 1;cactus_sprite[5][40][40] = 1;cactus_sprite[5][40][41] = 1;cactus_sprite[5][40][42] = 1;cactus_sprite[5][40][43] = 1;cactus_sprite[5][40][44] = 1;cactus_sprite[5][40][45] = 1;cactus_sprite[5][40][46] = 1;cactus_sprite[5][40][47] = 1;cactus_sprite[5][40][48] = 1;cactus_sprite[5][40][49] = 1;cactus_sprite[5][40][50] = 1;cactus_sprite[5][40][51] = 1;cactus_sprite[5][40][52] = 1;cactus_sprite[5][40][53] = 1;cactus_sprite[5][40][54] = 1;cactus_sprite[5][40][55] = 1;cactus_sprite[5][40][56] = 1;cactus_sprite[5][40][57] = 1;cactus_sprite[5][40][58] = 1;cactus_sprite[5][40][59] = 1;cactus_sprite[5][40][60] = 1;cactus_sprite[5][40][61] = 1;cactus_sprite[5][40][62] = 1;cactus_sprite[5][40][63] = 1;cactus_sprite[5][41][28] = 1;cactus_sprite[5][41][29] = 1;cactus_sprite[5][41][30] = 1;cactus_sprite[5][41][31] = 1;cactus_sprite[5][41][32] = 1;cactus_sprite[5][41][33] = 1;cactus_sprite[5][41][34] = 1;cactus_sprite[5][41][35] = 1;cactus_sprite[5][41][36] = 1;cactus_sprite[5][41][37] = 1;cactus_sprite[5][41][38] = 1;cactus_sprite[5][41][39] = 1;cactus_sprite[5][41][40] = 1;cactus_sprite[5][41][41] = 1;cactus_sprite[5][41][42] = 1;cactus_sprite[5][41][43] = 1;cactus_sprite[5][41][44] = 1;cactus_sprite[5][41][45] = 1;cactus_sprite[5][41][46] = 1;cactus_sprite[5][41][47] = 1;cactus_sprite[5][41][48] = 1;cactus_sprite[5][41][49] = 1;cactus_sprite[5][41][50] = 1;cactus_sprite[5][41][51] = 1;cactus_sprite[5][41][52] = 1;cactus_sprite[5][41][53] = 1;cactus_sprite[5][41][54] = 1;cactus_sprite[5][41][55] = 1;cactus_sprite[5][41][56] = 1;cactus_sprite[5][41][57] = 1;cactus_sprite[5][41][58] = 1;cactus_sprite[5][41][59] = 1;cactus_sprite[5][41][60] = 1;cactus_sprite[5][41][61] = 1;cactus_sprite[5][41][62] = 1;cactus_sprite[5][41][63] = 1;cactus_sprite[5][42][28] = 1;cactus_sprite[5][42][29] = 1;cactus_sprite[5][42][30] = 1;cactus_sprite[5][42][31] = 1;cactus_sprite[5][42][32] = 1;cactus_sprite[5][42][33] = 1;cactus_sprite[5][42][34] = 1;cactus_sprite[5][42][35] = 1;cactus_sprite[5][42][36] = 1;cactus_sprite[5][42][37] = 1;cactus_sprite[5][42][38] = 1;cactus_sprite[5][42][39] = 1;cactus_sprite[5][42][40] = 1;cactus_sprite[5][42][41] = 1;cactus_sprite[5][42][42] = 1;cactus_sprite[5][42][43] = 1;cactus_sprite[5][42][44] = 1;cactus_sprite[5][42][45] = 1;cactus_sprite[5][42][46] = 1;cactus_sprite[5][42][47] = 1;cactus_sprite[5][42][48] = 1;cactus_sprite[5][42][49] = 1;cactus_sprite[5][42][50] = 1;cactus_sprite[5][42][51] = 1;cactus_sprite[5][42][52] = 1;cactus_sprite[5][42][53] = 1;cactus_sprite[5][42][54] = 1;cactus_sprite[5][42][55] = 1;cactus_sprite[5][42][56] = 1;cactus_sprite[5][42][57] = 1;cactus_sprite[5][42][58] = 1;cactus_sprite[5][42][59] = 1;cactus_sprite[5][42][60] = 1;cactus_sprite[5][42][61] = 1;cactus_sprite[5][43][28] = 1;cactus_sprite[5][43][29] = 1;cactus_sprite[5][43][30] = 1;cactus_sprite[5][43][31] = 1;cactus_sprite[5][43][32] = 1;cactus_sprite[5][43][33] = 1;cactus_sprite[5][43][34] = 1;cactus_sprite[5][43][35] = 1;cactus_sprite[5][43][36] = 1;cactus_sprite[5][43][37] = 1;cactus_sprite[5][43][38] = 1;cactus_sprite[5][43][39] = 1;cactus_sprite[5][43][40] = 1;cactus_sprite[5][43][41] = 1;cactus_sprite[5][43][42] = 1;cactus_sprite[5][43][43] = 1;cactus_sprite[5][43][44] = 1;cactus_sprite[5][43][45] = 1;cactus_sprite[5][43][46] = 1;cactus_sprite[5][43][47] = 1;cactus_sprite[5][43][48] = 1;cactus_sprite[5][43][49] = 1;cactus_sprite[5][43][50] = 1;cactus_sprite[5][43][51] = 1;cactus_sprite[5][43][52] = 1;cactus_sprite[5][43][53] = 1;cactus_sprite[5][43][54] = 1;cactus_sprite[5][43][55] = 1;cactus_sprite[5][43][56] = 1;cactus_sprite[5][43][57] = 1;cactus_sprite[5][43][58] = 1;cactus_sprite[5][43][59] = 1;cactus_sprite[5][43][60] = 1;cactus_sprite[5][43][61] = 1;cactus_sprite[5][44][28] = 1;cactus_sprite[5][44][29] = 1;cactus_sprite[5][44][30] = 1;cactus_sprite[5][44][31] = 1;cactus_sprite[5][44][32] = 1;cactus_sprite[5][44][33] = 1;cactus_sprite[5][44][34] = 1;cactus_sprite[5][44][35] = 1;cactus_sprite[5][44][36] = 1;cactus_sprite[5][44][37] = 1;cactus_sprite[5][44][38] = 1;cactus_sprite[5][44][39] = 1;cactus_sprite[5][44][40] = 1;cactus_sprite[5][44][41] = 1;cactus_sprite[5][44][42] = 1;cactus_sprite[5][44][43] = 1;cactus_sprite[5][44][44] = 1;cactus_sprite[5][44][45] = 1;cactus_sprite[5][44][46] = 1;cactus_sprite[5][44][47] = 1;cactus_sprite[5][44][48] = 1;cactus_sprite[5][44][49] = 1;cactus_sprite[5][44][50] = 1;cactus_sprite[5][44][51] = 1;cactus_sprite[5][44][52] = 1;cactus_sprite[5][44][53] = 1;cactus_sprite[5][44][54] = 1;cactus_sprite[5][44][55] = 1;cactus_sprite[5][44][56] = 1;cactus_sprite[5][44][57] = 1;cactus_sprite[5][44][58] = 1;cactus_sprite[5][44][59] = 1;cactus_sprite[5][45][28] = 1;cactus_sprite[5][45][29] = 1;cactus_sprite[5][45][30] = 1;cactus_sprite[5][45][31] = 1;cactus_sprite[5][45][32] = 1;cactus_sprite[5][45][33] = 1;cactus_sprite[5][45][34] = 1;cactus_sprite[5][45][35] = 1;cactus_sprite[5][45][36] = 1;cactus_sprite[5][45][37] = 1;cactus_sprite[5][45][38] = 1;cactus_sprite[5][45][39] = 1;cactus_sprite[5][45][40] = 1;cactus_sprite[5][45][41] = 1;cactus_sprite[5][45][42] = 1;cactus_sprite[5][45][43] = 1;cactus_sprite[5][45][44] = 1;cactus_sprite[5][45][45] = 1;cactus_sprite[5][45][46] = 1;cactus_sprite[5][45][47] = 1;cactus_sprite[5][45][48] = 1;cactus_sprite[5][45][49] = 1;cactus_sprite[5][45][50] = 1;cactus_sprite[5][45][51] = 1;cactus_sprite[5][45][52] = 1;cactus_sprite[5][45][53] = 1;cactus_sprite[5][45][54] = 1;cactus_sprite[5][45][55] = 1;cactus_sprite[5][45][56] = 1;cactus_sprite[5][45][57] = 1;cactus_sprite[5][45][58] = 1;cactus_sprite[5][45][59] = 1;cactus_sprite[5][46][30] = 1;cactus_sprite[5][46][31] = 1;cactus_sprite[5][46][32] = 1;cactus_sprite[5][46][33] = 1;cactus_sprite[5][46][34] = 1;cactus_sprite[5][46][35] = 1;cactus_sprite[5][46][36] = 1;cactus_sprite[5][46][37] = 1;cactus_sprite[5][46][38] = 1;cactus_sprite[5][46][39] = 1;cactus_sprite[5][46][40] = 1;cactus_sprite[5][46][41] = 1;cactus_sprite[5][46][42] = 1;cactus_sprite[5][46][43] = 1;cactus_sprite[5][46][44] = 1;cactus_sprite[5][46][45] = 1;cactus_sprite[5][46][46] = 1;cactus_sprite[5][46][47] = 1;cactus_sprite[5][46][48] = 1;cactus_sprite[5][46][49] = 1;cactus_sprite[5][46][50] = 1;cactus_sprite[5][46][51] = 1;cactus_sprite[5][46][52] = 1;cactus_sprite[5][46][53] = 1;cactus_sprite[5][46][54] = 1;cactus_sprite[5][46][55] = 1;cactus_sprite[5][46][56] = 1;cactus_sprite[5][46][57] = 1;cactus_sprite[5][47][30] = 1;cactus_sprite[5][47][31] = 1;cactus_sprite[5][47][32] = 1;cactus_sprite[5][47][33] = 1;cactus_sprite[5][47][34] = 1;cactus_sprite[5][47][35] = 1;cactus_sprite[5][47][36] = 1;cactus_sprite[5][47][37] = 1;cactus_sprite[5][47][38] = 1;cactus_sprite[5][47][39] = 1;cactus_sprite[5][47][40] = 1;cactus_sprite[5][47][41] = 1;cactus_sprite[5][47][42] = 1;cactus_sprite[5][47][43] = 1;cactus_sprite[5][47][44] = 1;cactus_sprite[5][47][45] = 1;cactus_sprite[5][47][46] = 1;cactus_sprite[5][47][47] = 1;cactus_sprite[5][47][48] = 1;cactus_sprite[5][47][49] = 1;cactus_sprite[5][47][50] = 1;cactus_sprite[5][47][51] = 1;cactus_sprite[5][47][52] = 1;cactus_sprite[5][47][53] = 1;cactus_sprite[5][47][54] = 1;cactus_sprite[5][47][55] = 1;cactus_sprite[5][47][56] = 1;cactus_sprite[5][47][57] = 1;
	cactus_sprite[6][2][56] = 1;cactus_sprite[6][2][57] = 1;cactus_sprite[6][2][58] = 1;cactus_sprite[6][2][59] = 1;cactus_sprite[6][2][60] = 1;cactus_sprite[6][2][61] = 1;cactus_sprite[6][2][62] = 1;cactus_sprite[6][2][63] = 1;cactus_sprite[6][2][64] = 1;cactus_sprite[6][2][65] = 1;cactus_sprite[6][2][66] = 1;cactus_sprite[6][2][67] = 1;cactus_sprite[6][2][68] = 1;cactus_sprite[6][2][69] = 1;cactus_sprite[6][2][70] = 1;cactus_sprite[6][2][71] = 1;cactus_sprite[6][2][72] = 1;cactus_sprite[6][2][73] = 1;cactus_sprite[6][3][56] = 1;cactus_sprite[6][3][57] = 1;cactus_sprite[6][3][58] = 1;cactus_sprite[6][3][59] = 1;cactus_sprite[6][3][60] = 1;cactus_sprite[6][3][61] = 1;cactus_sprite[6][3][62] = 1;cactus_sprite[6][3][63] = 1;cactus_sprite[6][3][64] = 1;cactus_sprite[6][3][65] = 1;cactus_sprite[6][3][66] = 1;cactus_sprite[6][3][67] = 1;cactus_sprite[6][3][68] = 1;cactus_sprite[6][3][69] = 1;cactus_sprite[6][3][70] = 1;cactus_sprite[6][3][71] = 1;cactus_sprite[6][3][72] = 1;cactus_sprite[6][3][73] = 1;cactus_sprite[6][4][54] = 1;cactus_sprite[6][4][55] = 1;cactus_sprite[6][4][56] = 1;cactus_sprite[6][4][57] = 1;cactus_sprite[6][4][58] = 1;cactus_sprite[6][4][59] = 1;cactus_sprite[6][4][60] = 1;cactus_sprite[6][4][61] = 1;cactus_sprite[6][4][62] = 1;cactus_sprite[6][4][63] = 1;cactus_sprite[6][4][64] = 1;cactus_sprite[6][4][65] = 1;cactus_sprite[6][4][66] = 1;cactus_sprite[6][4][67] = 1;cactus_sprite[6][4][68] = 1;cactus_sprite[6][4][69] = 1;cactus_sprite[6][4][70] = 1;cactus_sprite[6][4][71] = 1;cactus_sprite[6][4][72] = 1;cactus_sprite[6][4][73] = 1;cactus_sprite[6][4][74] = 1;cactus_sprite[6][4][75] = 1;cactus_sprite[6][5][54] = 1;cactus_sprite[6][5][55] = 1;cactus_sprite[6][5][56] = 1;cactus_sprite[6][5][57] = 1;cactus_sprite[6][5][58] = 1;cactus_sprite[6][5][59] = 1;cactus_sprite[6][5][60] = 1;cactus_sprite[6][5][61] = 1;cactus_sprite[6][5][62] = 1;cactus_sprite[6][5][63] = 1;cactus_sprite[6][5][64] = 1;cactus_sprite[6][5][65] = 1;cactus_sprite[6][5][66] = 1;cactus_sprite[6][5][67] = 1;cactus_sprite[6][5][68] = 1;cactus_sprite[6][5][69] = 1;cactus_sprite[6][5][70] = 1;cactus_sprite[6][5][71] = 1;cactus_sprite[6][5][72] = 1;cactus_sprite[6][5][73] = 1;cactus_sprite[6][5][74] = 1;cactus_sprite[6][5][75] = 1;cactus_sprite[6][6][56] = 1;cactus_sprite[6][6][57] = 1;cactus_sprite[6][6][58] = 1;cactus_sprite[6][6][59] = 1;cactus_sprite[6][6][60] = 1;cactus_sprite[6][6][61] = 1;cactus_sprite[6][6][62] = 1;cactus_sprite[6][6][63] = 1;cactus_sprite[6][6][64] = 1;cactus_sprite[6][6][65] = 1;cactus_sprite[6][6][66] = 1;cactus_sprite[6][6][67] = 1;cactus_sprite[6][6][68] = 1;cactus_sprite[6][6][69] = 1;cactus_sprite[6][6][70] = 1;cactus_sprite[6][6][71] = 1;cactus_sprite[6][6][72] = 1;cactus_sprite[6][6][73] = 1;cactus_sprite[6][6][74] = 1;cactus_sprite[6][6][75] = 1;cactus_sprite[6][6][76] = 1;cactus_sprite[6][6][77] = 1;cactus_sprite[6][7][56] = 1;cactus_sprite[6][7][57] = 1;cactus_sprite[6][7][58] = 1;cactus_sprite[6][7][59] = 1;cactus_sprite[6][7][60] = 1;cactus_sprite[6][7][61] = 1;cactus_sprite[6][7][62] = 1;cactus_sprite[6][7][63] = 1;cactus_sprite[6][7][64] = 1;cactus_sprite[6][7][65] = 1;cactus_sprite[6][7][66] = 1;cactus_sprite[6][7][67] = 1;cactus_sprite[6][7][68] = 1;cactus_sprite[6][7][69] = 1;cactus_sprite[6][7][70] = 1;cactus_sprite[6][7][71] = 1;cactus_sprite[6][7][72] = 1;cactus_sprite[6][7][73] = 1;cactus_sprite[6][7][74] = 1;cactus_sprite[6][7][75] = 1;cactus_sprite[6][7][76] = 1;cactus_sprite[6][7][77] = 1;cactus_sprite[6][8][74] = 1;cactus_sprite[6][8][75] = 1;cactus_sprite[6][8][76] = 1;cactus_sprite[6][8][77] = 1;cactus_sprite[6][8][78] = 1;cactus_sprite[6][8][79] = 1;cactus_sprite[6][9][74] = 1;cactus_sprite[6][9][75] = 1;cactus_sprite[6][9][76] = 1;cactus_sprite[6][9][77] = 1;cactus_sprite[6][9][78] = 1;cactus_sprite[6][9][79] = 1;cactus_sprite[6][10][74] = 1;cactus_sprite[6][10][75] = 1;cactus_sprite[6][10][76] = 1;cactus_sprite[6][10][77] = 1;cactus_sprite[6][10][78] = 1;cactus_sprite[6][10][79] = 1;cactus_sprite[6][11][74] = 1;cactus_sprite[6][11][75] = 1;cactus_sprite[6][11][76] = 1;cactus_sprite[6][11][77] = 1;cactus_sprite[6][11][78] = 1;cactus_sprite[6][11][79] = 1;cactus_sprite[6][12][46] = 1;cactus_sprite[6][12][47] = 1;cactus_sprite[6][12][48] = 1;cactus_sprite[6][12][49] = 1;cactus_sprite[6][12][50] = 1;cactus_sprite[6][12][51] = 1;cactus_sprite[6][12][52] = 1;cactus_sprite[6][12][53] = 1;cactus_sprite[6][12][54] = 1;cactus_sprite[6][12][55] = 1;cactus_sprite[6][12][56] = 1;cactus_sprite[6][12][57] = 1;cactus_sprite[6][12][58] = 1;cactus_sprite[6][12][59] = 1;cactus_sprite[6][12][60] = 1;cactus_sprite[6][12][61] = 1;cactus_sprite[6][12][62] = 1;cactus_sprite[6][12][63] = 1;cactus_sprite[6][12][64] = 1;cactus_sprite[6][12][65] = 1;cactus_sprite[6][12][66] = 1;cactus_sprite[6][12][67] = 1;cactus_sprite[6][12][68] = 1;cactus_sprite[6][12][69] = 1;cactus_sprite[6][12][70] = 1;cactus_sprite[6][12][71] = 1;cactus_sprite[6][12][72] = 1;cactus_sprite[6][12][73] = 1;cactus_sprite[6][12][74] = 1;cactus_sprite[6][12][75] = 1;cactus_sprite[6][12][76] = 1;cactus_sprite[6][12][77] = 1;cactus_sprite[6][12][78] = 1;cactus_sprite[6][12][79] = 1;cactus_sprite[6][12][80] = 1;cactus_sprite[6][12][81] = 1;cactus_sprite[6][12][82] = 1;cactus_sprite[6][12][83] = 1;cactus_sprite[6][12][84] = 1;cactus_sprite[6][12][85] = 1;cactus_sprite[6][12][86] = 1;cactus_sprite[6][12][87] = 1;cactus_sprite[6][12][88] = 1;cactus_sprite[6][12][89] = 1;cactus_sprite[6][12][90] = 1;cactus_sprite[6][12][91] = 1;cactus_sprite[6][12][92] = 1;cactus_sprite[6][12][93] = 1;cactus_sprite[6][12][94] = 1;cactus_sprite[6][12][95] = 1;cactus_sprite[6][12][96] = 1;cactus_sprite[6][12][97] = 1;cactus_sprite[6][12][98] = 1;cactus_sprite[6][12][99] = 1;cactus_sprite[6][13][46] = 1;cactus_sprite[6][13][47] = 1;cactus_sprite[6][13][48] = 1;cactus_sprite[6][13][49] = 1;cactus_sprite[6][13][50] = 1;cactus_sprite[6][13][51] = 1;cactus_sprite[6][13][52] = 1;cactus_sprite[6][13][53] = 1;cactus_sprite[6][13][54] = 1;cactus_sprite[6][13][55] = 1;cactus_sprite[6][13][56] = 1;cactus_sprite[6][13][57] = 1;cactus_sprite[6][13][58] = 1;cactus_sprite[6][13][59] = 1;cactus_sprite[6][13][60] = 1;cactus_sprite[6][13][61] = 1;cactus_sprite[6][13][62] = 1;cactus_sprite[6][13][63] = 1;cactus_sprite[6][13][64] = 1;cactus_sprite[6][13][65] = 1;cactus_sprite[6][13][66] = 1;cactus_sprite[6][13][67] = 1;cactus_sprite[6][13][68] = 1;cactus_sprite[6][13][69] = 1;cactus_sprite[6][13][70] = 1;cactus_sprite[6][13][71] = 1;cactus_sprite[6][13][72] = 1;cactus_sprite[6][13][73] = 1;cactus_sprite[6][13][74] = 1;cactus_sprite[6][13][75] = 1;cactus_sprite[6][13][76] = 1;cactus_sprite[6][13][77] = 1;cactus_sprite[6][13][78] = 1;cactus_sprite[6][13][79] = 1;cactus_sprite[6][13][80] = 1;cactus_sprite[6][13][81] = 1;cactus_sprite[6][13][82] = 1;cactus_sprite[6][13][83] = 1;cactus_sprite[6][13][84] = 1;cactus_sprite[6][13][85] = 1;cactus_sprite[6][13][86] = 1;cactus_sprite[6][13][87] = 1;cactus_sprite[6][13][88] = 1;cactus_sprite[6][13][89] = 1;cactus_sprite[6][13][90] = 1;cactus_sprite[6][13][91] = 1;cactus_sprite[6][13][92] = 1;cactus_sprite[6][13][93] = 1;cactus_sprite[6][13][94] = 1;cactus_sprite[6][13][95] = 1;cactus_sprite[6][13][96] = 1;cactus_sprite[6][13][97] = 1;cactus_sprite[6][13][98] = 1;cactus_sprite[6][13][99] = 1;cactus_sprite[6][14][44] = 1;cactus_sprite[6][14][45] = 1;cactus_sprite[6][14][46] = 1;cactus_sprite[6][14][47] = 1;cactus_sprite[6][14][48] = 1;cactus_sprite[6][14][49] = 1;cactus_sprite[6][14][50] = 1;cactus_sprite[6][14][51] = 1;cactus_sprite[6][14][52] = 1;cactus_sprite[6][14][53] = 1;cactus_sprite[6][14][54] = 1;cactus_sprite[6][14][55] = 1;cactus_sprite[6][14][56] = 1;cactus_sprite[6][14][57] = 1;cactus_sprite[6][14][58] = 1;cactus_sprite[6][14][59] = 1;cactus_sprite[6][14][60] = 1;cactus_sprite[6][14][61] = 1;cactus_sprite[6][14][62] = 1;cactus_sprite[6][14][63] = 1;cactus_sprite[6][14][64] = 1;cactus_sprite[6][14][65] = 1;cactus_sprite[6][14][66] = 1;cactus_sprite[6][14][67] = 1;cactus_sprite[6][14][68] = 1;cactus_sprite[6][14][69] = 1;cactus_sprite[6][14][70] = 1;cactus_sprite[6][14][71] = 1;cactus_sprite[6][14][72] = 1;cactus_sprite[6][14][73] = 1;cactus_sprite[6][14][74] = 1;cactus_sprite[6][14][75] = 1;cactus_sprite[6][14][76] = 1;cactus_sprite[6][14][77] = 1;cactus_sprite[6][14][78] = 1;cactus_sprite[6][14][79] = 1;cactus_sprite[6][14][80] = 1;cactus_sprite[6][14][81] = 1;cactus_sprite[6][14][82] = 1;cactus_sprite[6][14][83] = 1;cactus_sprite[6][14][84] = 1;cactus_sprite[6][14][85] = 1;cactus_sprite[6][14][86] = 1;cactus_sprite[6][14][87] = 1;cactus_sprite[6][14][88] = 1;cactus_sprite[6][14][89] = 1;cactus_sprite[6][14][90] = 1;cactus_sprite[6][14][91] = 1;cactus_sprite[6][14][92] = 1;cactus_sprite[6][14][93] = 1;cactus_sprite[6][14][94] = 1;cactus_sprite[6][14][95] = 1;cactus_sprite[6][14][96] = 1;cactus_sprite[6][14][97] = 1;cactus_sprite[6][14][98] = 1;cactus_sprite[6][14][99] = 1;cactus_sprite[6][15][44] = 1;cactus_sprite[6][15][45] = 1;cactus_sprite[6][15][46] = 1;cactus_sprite[6][15][47] = 1;cactus_sprite[6][15][48] = 1;cactus_sprite[6][15][49] = 1;cactus_sprite[6][15][50] = 1;cactus_sprite[6][15][51] = 1;cactus_sprite[6][15][52] = 1;cactus_sprite[6][15][53] = 1;cactus_sprite[6][15][54] = 1;cactus_sprite[6][15][55] = 1;cactus_sprite[6][15][56] = 1;cactus_sprite[6][15][57] = 1;cactus_sprite[6][15][58] = 1;cactus_sprite[6][15][59] = 1;cactus_sprite[6][15][60] = 1;cactus_sprite[6][15][61] = 1;cactus_sprite[6][15][62] = 1;cactus_sprite[6][15][63] = 1;cactus_sprite[6][15][64] = 1;cactus_sprite[6][15][65] = 1;cactus_sprite[6][15][66] = 1;cactus_sprite[6][15][67] = 1;cactus_sprite[6][15][68] = 1;cactus_sprite[6][15][69] = 1;cactus_sprite[6][15][70] = 1;cactus_sprite[6][15][71] = 1;cactus_sprite[6][15][72] = 1;cactus_sprite[6][15][73] = 1;cactus_sprite[6][15][74] = 1;cactus_sprite[6][15][75] = 1;cactus_sprite[6][15][76] = 1;cactus_sprite[6][15][77] = 1;cactus_sprite[6][15][78] = 1;cactus_sprite[6][15][79] = 1;cactus_sprite[6][15][80] = 1;cactus_sprite[6][15][81] = 1;cactus_sprite[6][15][82] = 1;cactus_sprite[6][15][83] = 1;cactus_sprite[6][15][84] = 1;cactus_sprite[6][15][85] = 1;cactus_sprite[6][15][86] = 1;cactus_sprite[6][15][87] = 1;cactus_sprite[6][15][88] = 1;cactus_sprite[6][15][89] = 1;cactus_sprite[6][15][90] = 1;cactus_sprite[6][15][91] = 1;cactus_sprite[6][15][92] = 1;cactus_sprite[6][15][93] = 1;cactus_sprite[6][15][94] = 1;cactus_sprite[6][15][95] = 1;cactus_sprite[6][15][96] = 1;cactus_sprite[6][15][97] = 1;cactus_sprite[6][15][98] = 1;cactus_sprite[6][15][99] = 1;cactus_sprite[6][16][46] = 1;cactus_sprite[6][16][47] = 1;cactus_sprite[6][16][48] = 1;cactus_sprite[6][16][49] = 1;cactus_sprite[6][16][50] = 1;cactus_sprite[6][16][51] = 1;cactus_sprite[6][16][52] = 1;cactus_sprite[6][16][53] = 1;cactus_sprite[6][16][54] = 1;cactus_sprite[6][16][55] = 1;cactus_sprite[6][16][56] = 1;cactus_sprite[6][16][57] = 1;cactus_sprite[6][16][58] = 1;cactus_sprite[6][16][59] = 1;cactus_sprite[6][16][60] = 1;cactus_sprite[6][16][61] = 1;cactus_sprite[6][16][62] = 1;cactus_sprite[6][16][63] = 1;cactus_sprite[6][16][64] = 1;cactus_sprite[6][16][65] = 1;cactus_sprite[6][16][66] = 1;cactus_sprite[6][16][67] = 1;cactus_sprite[6][16][68] = 1;cactus_sprite[6][16][69] = 1;cactus_sprite[6][16][70] = 1;cactus_sprite[6][16][71] = 1;cactus_sprite[6][16][72] = 1;cactus_sprite[6][16][73] = 1;cactus_sprite[6][16][74] = 1;cactus_sprite[6][16][75] = 1;cactus_sprite[6][16][76] = 1;cactus_sprite[6][16][77] = 1;cactus_sprite[6][16][78] = 1;cactus_sprite[6][16][79] = 1;cactus_sprite[6][16][80] = 1;cactus_sprite[6][16][81] = 1;cactus_sprite[6][16][82] = 1;cactus_sprite[6][16][83] = 1;cactus_sprite[6][16][84] = 1;cactus_sprite[6][16][85] = 1;cactus_sprite[6][16][86] = 1;cactus_sprite[6][16][87] = 1;cactus_sprite[6][16][88] = 1;cactus_sprite[6][16][89] = 1;cactus_sprite[6][16][90] = 1;cactus_sprite[6][16][91] = 1;cactus_sprite[6][16][92] = 1;cactus_sprite[6][16][93] = 1;cactus_sprite[6][16][94] = 1;cactus_sprite[6][16][95] = 1;cactus_sprite[6][16][96] = 1;cactus_sprite[6][16][97] = 1;cactus_sprite[6][16][98] = 1;cactus_sprite[6][16][99] = 1;cactus_sprite[6][17][46] = 1;cactus_sprite[6][17][47] = 1;cactus_sprite[6][17][48] = 1;cactus_sprite[6][17][49] = 1;cactus_sprite[6][17][50] = 1;cactus_sprite[6][17][51] = 1;cactus_sprite[6][17][52] = 1;cactus_sprite[6][17][53] = 1;cactus_sprite[6][17][54] = 1;cactus_sprite[6][17][55] = 1;cactus_sprite[6][17][56] = 1;cactus_sprite[6][17][57] = 1;cactus_sprite[6][17][58] = 1;cactus_sprite[6][17][59] = 1;cactus_sprite[6][17][60] = 1;cactus_sprite[6][17][61] = 1;cactus_sprite[6][17][62] = 1;cactus_sprite[6][17][63] = 1;cactus_sprite[6][17][64] = 1;cactus_sprite[6][17][65] = 1;cactus_sprite[6][17][66] = 1;cactus_sprite[6][17][67] = 1;cactus_sprite[6][17][68] = 1;cactus_sprite[6][17][69] = 1;cactus_sprite[6][17][70] = 1;cactus_sprite[6][17][71] = 1;cactus_sprite[6][17][72] = 1;cactus_sprite[6][17][73] = 1;cactus_sprite[6][17][74] = 1;cactus_sprite[6][17][75] = 1;cactus_sprite[6][17][76] = 1;cactus_sprite[6][17][77] = 1;cactus_sprite[6][17][78] = 1;cactus_sprite[6][17][79] = 1;cactus_sprite[6][17][80] = 1;cactus_sprite[6][17][81] = 1;cactus_sprite[6][17][82] = 1;cactus_sprite[6][17][83] = 1;cactus_sprite[6][17][84] = 1;cactus_sprite[6][17][85] = 1;cactus_sprite[6][17][86] = 1;cactus_sprite[6][17][87] = 1;cactus_sprite[6][17][88] = 1;cactus_sprite[6][17][89] = 1;cactus_sprite[6][17][90] = 1;cactus_sprite[6][17][91] = 1;cactus_sprite[6][17][92] = 1;cactus_sprite[6][17][93] = 1;cactus_sprite[6][17][94] = 1;cactus_sprite[6][17][95] = 1;cactus_sprite[6][17][96] = 1;cactus_sprite[6][17][97] = 1;cactus_sprite[6][17][98] = 1;cactus_sprite[6][17][99] = 1;cactus_sprite[6][18][74] = 1;cactus_sprite[6][18][75] = 1;cactus_sprite[6][18][76] = 1;cactus_sprite[6][18][77] = 1;cactus_sprite[6][19][74] = 1;cactus_sprite[6][19][75] = 1;cactus_sprite[6][19][76] = 1;cactus_sprite[6][19][77] = 1;cactus_sprite[6][20][74] = 1;cactus_sprite[6][20][75] = 1;cactus_sprite[6][20][76] = 1;cactus_sprite[6][20][77] = 1;cactus_sprite[6][21][74] = 1;cactus_sprite[6][21][75] = 1;cactus_sprite[6][21][76] = 1;cactus_sprite[6][21][77] = 1;cactus_sprite[6][22][56] = 1;cactus_sprite[6][22][57] = 1;cactus_sprite[6][22][58] = 1;cactus_sprite[6][22][59] = 1;cactus_sprite[6][22][60] = 1;cactus_sprite[6][22][61] = 1;cactus_sprite[6][22][62] = 1;cactus_sprite[6][22][63] = 1;cactus_sprite[6][22][64] = 1;cactus_sprite[6][22][65] = 1;cactus_sprite[6][22][66] = 1;cactus_sprite[6][22][67] = 1;cactus_sprite[6][22][68] = 1;cactus_sprite[6][22][69] = 1;cactus_sprite[6][22][70] = 1;cactus_sprite[6][22][71] = 1;cactus_sprite[6][22][72] = 1;cactus_sprite[6][22][73] = 1;cactus_sprite[6][22][74] = 1;cactus_sprite[6][22][75] = 1;cactus_sprite[6][22][76] = 1;cactus_sprite[6][22][77] = 1;cactus_sprite[6][23][56] = 1;cactus_sprite[6][23][57] = 1;cactus_sprite[6][23][58] = 1;cactus_sprite[6][23][59] = 1;cactus_sprite[6][23][60] = 1;cactus_sprite[6][23][61] = 1;cactus_sprite[6][23][62] = 1;cactus_sprite[6][23][63] = 1;cactus_sprite[6][23][64] = 1;cactus_sprite[6][23][65] = 1;cactus_sprite[6][23][66] = 1;cactus_sprite[6][23][67] = 1;cactus_sprite[6][23][68] = 1;cactus_sprite[6][23][69] = 1;cactus_sprite[6][23][70] = 1;cactus_sprite[6][23][71] = 1;cactus_sprite[6][23][72] = 1;cactus_sprite[6][23][73] = 1;cactus_sprite[6][23][74] = 1;cactus_sprite[6][23][75] = 1;cactus_sprite[6][23][76] = 1;cactus_sprite[6][23][77] = 1;cactus_sprite[6][24][54] = 1;cactus_sprite[6][24][55] = 1;cactus_sprite[6][24][56] = 1;cactus_sprite[6][24][57] = 1;cactus_sprite[6][24][58] = 1;cactus_sprite[6][24][59] = 1;cactus_sprite[6][24][60] = 1;cactus_sprite[6][24][61] = 1;cactus_sprite[6][24][62] = 1;cactus_sprite[6][24][63] = 1;cactus_sprite[6][24][64] = 1;cactus_sprite[6][24][65] = 1;cactus_sprite[6][24][66] = 1;cactus_sprite[6][24][67] = 1;cactus_sprite[6][24][68] = 1;cactus_sprite[6][24][69] = 1;cactus_sprite[6][24][70] = 1;cactus_sprite[6][24][71] = 1;cactus_sprite[6][24][72] = 1;cactus_sprite[6][24][73] = 1;cactus_sprite[6][24][74] = 1;cactus_sprite[6][24][75] = 1;cactus_sprite[6][25][54] = 1;cactus_sprite[6][25][55] = 1;cactus_sprite[6][25][56] = 1;cactus_sprite[6][25][57] = 1;cactus_sprite[6][25][58] = 1;cactus_sprite[6][25][59] = 1;cactus_sprite[6][25][60] = 1;cactus_sprite[6][25][61] = 1;cactus_sprite[6][25][62] = 1;cactus_sprite[6][25][63] = 1;cactus_sprite[6][25][64] = 1;cactus_sprite[6][25][65] = 1;cactus_sprite[6][25][66] = 1;cactus_sprite[6][25][67] = 1;cactus_sprite[6][25][68] = 1;cactus_sprite[6][25][69] = 1;cactus_sprite[6][25][70] = 1;cactus_sprite[6][25][71] = 1;cactus_sprite[6][25][72] = 1;cactus_sprite[6][25][73] = 1;cactus_sprite[6][25][74] = 1;cactus_sprite[6][25][75] = 1;cactus_sprite[6][26][56] = 1;cactus_sprite[6][26][57] = 1;cactus_sprite[6][26][58] = 1;cactus_sprite[6][26][59] = 1;cactus_sprite[6][26][60] = 1;cactus_sprite[6][26][61] = 1;cactus_sprite[6][26][62] = 1;cactus_sprite[6][26][63] = 1;cactus_sprite[6][26][64] = 1;cactus_sprite[6][26][65] = 1;cactus_sprite[6][26][66] = 1;cactus_sprite[6][26][67] = 1;cactus_sprite[6][26][68] = 1;cactus_sprite[6][26][69] = 1;cactus_sprite[6][26][70] = 1;cactus_sprite[6][26][71] = 1;cactus_sprite[6][26][72] = 1;cactus_sprite[6][26][73] = 1;cactus_sprite[6][27][56] = 1;cactus_sprite[6][27][57] = 1;cactus_sprite[6][27][58] = 1;cactus_sprite[6][27][59] = 1;cactus_sprite[6][27][60] = 1;cactus_sprite[6][27][61] = 1;cactus_sprite[6][27][62] = 1;cactus_sprite[6][27][63] = 1;cactus_sprite[6][27][64] = 1;cactus_sprite[6][27][65] = 1;cactus_sprite[6][27][66] = 1;cactus_sprite[6][27][67] = 1;cactus_sprite[6][27][68] = 1;cactus_sprite[6][27][69] = 1;cactus_sprite[6][27][70] = 1;cactus_sprite[6][27][71] = 1;cactus_sprite[6][27][72] = 1;cactus_sprite[6][27][73] = 1;
	
	
	
	for(i=0; i < 4; i=i+1) begin
		cactus_x = count_h - (1024 - cactuses[i]);
		cactus_y = 100 - (ground_y - count_v);
		
		if(cactuses[i] == 0)
			choice = choice + 1;
		
		if ((cactus_x >= 0 && cactus_x < 50) && (cactus_y >= 0 && cactus_y < 100)) begin
			if (cactus_sprite[cactuses_sprite_choice[choice]][cactus_x][cactus_y] == 1) begin
				r = 1;
				g = 1;
				b = 1;
			end
		end
	end
	
	// -- FRAME --
	if(count_v < 6 & count_v >= 0) begin r = 1;g = 1;b = 1; end
	if(count_v <= 768 & count_v > 768 - 5) begin r = 1;g = 1;b = 1; end
	if(count_h <= 1024 & count_h > 1024 - 6) begin r = 1;g = 1;b = 1; end
	if(count_h > 0 & count_h <= 5) begin r = 1;g = 1;b = 1; end
	// --
end
else begin
	r = 0;
	g = 0;
	b = 0;
end
end
endmodule
